//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Wed Jan 31 16:31:54 2024
// Version: 2023.2 2023.2.0.10
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// BVF_RISCV_SUBSYSTEM
module BVF_RISCV_SUBSYSTEM(
    // Inputs
    ADC_IRQn,
    CAPE_APB_MTARGET_PRDATAS1,
    CAPE_APB_MTARGET_PREADYS1,
    CAPE_APB_MTARGET_PSLVERRS1,
    CSI_APB_MTARGET_PRDATAS2,
    CSI_APB_MTARGET_PREADYS2,
    CSI_APB_MTARGET_PSLVERRS2,
    EMMC_STRB,
    FIC_0_ACLK,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARREADY,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWREADY,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BRESP,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BVALID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RDATA,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RLAST,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RRESP,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RVALID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WREADY,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARADDR,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARBURST,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARCACHE,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLEN,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLOCK,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARPROT,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARQOS,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARSIZE,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARVALID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWADDR,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWBURST,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWCACHE,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLEN,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLOCK,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWPROT,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWQOS,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWSIZE,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWVALID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BREADY,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RREADY,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WDATA,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WLAST,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WSTRB,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WVALID,
    FIC_1_ACLK,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARREADY,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWREADY,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BRESP,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BVALID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RDATA,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RLAST,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RRESP,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RVALID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WREADY,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARADDR,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARBURST,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARCACHE,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLEN,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLOCK,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARPROT,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARQOS,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARSIZE,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARVALID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWADDR,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWBURST,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWCACHE,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLEN,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLOCK,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWPROT,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWQOS,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWSIZE,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWVALID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BREADY,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RREADY,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WDATA,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WLAST,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WSTRB,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WVALID,
    FIC_2_ACLK,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARADDR,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARBURST,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARCACHE,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLEN,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLOCK,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARPROT,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARQOS,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARSIZE,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARVALID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWADDR,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWBURST,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWCACHE,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLEN,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLOCK,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWPROT,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWQOS,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWSIZE,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWVALID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BREADY,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RREADY,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WDATA,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WLAST,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WSTRB,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WVALID,
    FIC_3_PCLK,
    GPIO_2_F2M,
    HSI_APB_MTARGET_PRDATAS4,
    HSI_APB_MTARGET_PREADYS4,
    HSI_APB_MTARGET_PSLVERRS4,
    M2_APB_MTARGET_PRDATAS16,
    M2_APB_MTARGET_PREADYS16,
    M2_APB_MTARGET_PSLVERRS16,
    M2_UART_CTS,
    M2_UART_RXD,
    MAC_1_MDI_F2M,
    MMUART_2_RXD,
    MMUART_3_RXD,
    MMUART_4_RXD,
    MSS_INT_F2M,
    PCIE_INT,
    PHY_INTn,
    PRESETN,
    REFCLK,
    REFCLK_N,
    SD_DET,
    SGMII_RX0_N,
    SGMII_RX0_P,
    SGMII_RX1_N,
    SGMII_RX1_P,
    SPI_0_DI,
    SPI_1_DI,
    UART0_RXD,
    USB_CLK,
    USB_DIR,
    USB_NXT,
    USB_OCn,
    USER_BUTTON,
    // Outputs
    ADC_CSn,
    ADC_SCK,
    CA,
    CAPE_APB_MTARGET_PADDRS,
    CAPE_APB_MTARGET_PENABLES,
    CAPE_APB_MTARGET_PSELS1,
    CAPE_APB_MTARGET_PWDATAS,
    CAPE_APB_MTARGET_PWRITES,
    CK,
    CKE,
    CK_N,
    CS,
    CSI_APB_MTARGET_PSELS2,
    DM,
    EMMC_CLK,
    EMMC_RSTN,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARADDR,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARBURST,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARCACHE,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARLEN,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARLOCK,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARPROT,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARQOS,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARSIZE,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARVALID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWADDR,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWBURST,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWCACHE,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWLEN,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWLOCK,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWPROT,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWQOS,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWSIZE,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWVALID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BREADY,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RREADY,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WDATA,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WLAST,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WSTRB,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WVALID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARREADY,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWREADY,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BRESP,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BVALID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RDATA,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RLAST,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RRESP,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RVALID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WREADY,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARADDR,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARBURST,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARCACHE,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARLEN,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARLOCK,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARPROT,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARQOS,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARSIZE,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARVALID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWADDR,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWBURST,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWCACHE,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWLEN,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWLOCK,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWPROT,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWQOS,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWSIZE,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWVALID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BREADY,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RREADY,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WDATA,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WLAST,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WSTRB,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WVALID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARREADY,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWREADY,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BRESP,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BVALID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RDATA,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RLAST,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RRESP,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RVALID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WREADY,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARREADY,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWREADY,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BRESP,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BVALID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RDATA,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RLAST,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RRESP,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RVALID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WREADY,
    FIC_3_APB_M_PSTRB,
    GPIO_2_M2F,
    GPIO_2_OE_M2F,
    HSI_APB_MTARGET_PSELS4,
    M2_APB_MTARGET_PSELS16,
    M2_UART_RTS,
    M2_UART_TXD,
    M2_W_DISABLE1,
    M2_W_DISABLE2,
    MAC_1_MDC_M2F,
    MAC_1_MDO_M2F,
    MAC_1_MDO_OE_M2F,
    MMUART_2_TXD,
    MMUART_3_TXD,
    MMUART_4_TXD,
    MSS_DLL_LOCKS,
    MSS_RESET_N_M2F,
    ODT,
    PHY_MDC,
    RESET_N,
    SD_CARD_CS,
    SGMII_TX0_N,
    SGMII_TX0_P,
    SGMII_TX1_N,
    SGMII_TX1_P,
    SPI_0_CLK,
    SPI_0_DO,
    SPI_0_SS1,
    SPI_1_CLK,
    SPI_1_DO,
    SPI_1_SS1,
    UART0_TXD,
    USB_STP,
    VIO_ENABLE,
    // Inouts
    ADC_MISO,
    ADC_MOSI,
    DQ,
    DQS,
    DQS_N,
    EMMC_CMD,
    EMMC_DATA0,
    EMMC_DATA1,
    EMMC_DATA2,
    EMMC_DATA3,
    EMMC_DATA4,
    EMMC_DATA5,
    EMMC_DATA6,
    EMMC_DATA7,
    I2C0_SCL,
    I2C0_SDA,
    I2C_1_SCL,
    I2C_1_SDA,
    PHY_MDIO,
    USB_DATA0,
    USB_DATA1,
    USB_DATA2,
    USB_DATA3,
    USB_DATA4,
    USB_DATA5,
    USB_DATA6,
    USB_DATA7
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input         ADC_IRQn;
input  [31:0] CAPE_APB_MTARGET_PRDATAS1;
input         CAPE_APB_MTARGET_PREADYS1;
input         CAPE_APB_MTARGET_PSLVERRS1;
input  [31:0] CSI_APB_MTARGET_PRDATAS2;
input         CSI_APB_MTARGET_PREADYS2;
input         CSI_APB_MTARGET_PSLVERRS2;
input         EMMC_STRB;
input         FIC_0_ACLK;
input         FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARREADY;
input         FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWREADY;
input  [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BID;
input  [1:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BRESP;
input         FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BVALID;
input  [63:0] FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RDATA;
input  [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RID;
input         FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RLAST;
input  [1:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RRESP;
input         FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RVALID;
input         FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WREADY;
input  [37:0] FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARADDR;
input  [1:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARBURST;
input  [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARCACHE;
input  [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARID;
input  [7:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLEN;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLOCK;
input  [2:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARPROT;
input  [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARQOS;
input  [2:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARSIZE;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARVALID;
input  [37:0] FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWADDR;
input  [1:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWBURST;
input  [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWCACHE;
input  [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWID;
input  [7:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLEN;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLOCK;
input  [2:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWPROT;
input  [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWQOS;
input  [2:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWSIZE;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWVALID;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BREADY;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RREADY;
input  [63:0] FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WDATA;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WLAST;
input  [7:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WSTRB;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WVALID;
input         FIC_1_ACLK;
input         FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARREADY;
input         FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWREADY;
input  [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BID;
input  [1:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BRESP;
input         FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BVALID;
input  [63:0] FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RDATA;
input  [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RID;
input         FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RLAST;
input  [1:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RRESP;
input         FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RVALID;
input         FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WREADY;
input  [37:0] FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARADDR;
input  [1:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARBURST;
input  [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARCACHE;
input  [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARID;
input  [7:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLEN;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLOCK;
input  [2:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARPROT;
input  [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARQOS;
input  [2:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARSIZE;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARVALID;
input  [37:0] FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWADDR;
input  [1:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWBURST;
input  [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWCACHE;
input  [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWID;
input  [7:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLEN;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLOCK;
input  [2:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWPROT;
input  [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWQOS;
input  [2:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWSIZE;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWVALID;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BREADY;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RREADY;
input  [63:0] FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WDATA;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WLAST;
input  [7:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WSTRB;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WVALID;
input         FIC_2_ACLK;
input  [37:0] FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARADDR;
input  [1:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARBURST;
input  [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARCACHE;
input  [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARID;
input  [7:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLEN;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLOCK;
input  [2:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARPROT;
input  [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARQOS;
input  [2:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARSIZE;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARVALID;
input  [37:0] FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWADDR;
input  [1:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWBURST;
input  [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWCACHE;
input  [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWID;
input  [7:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLEN;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLOCK;
input  [2:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWPROT;
input  [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWQOS;
input  [2:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWSIZE;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWVALID;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BREADY;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RREADY;
input  [63:0] FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WDATA;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WLAST;
input  [7:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WSTRB;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WVALID;
input         FIC_3_PCLK;
input  [27:0] GPIO_2_F2M;
input  [31:0] HSI_APB_MTARGET_PRDATAS4;
input         HSI_APB_MTARGET_PREADYS4;
input         HSI_APB_MTARGET_PSLVERRS4;
input  [31:0] M2_APB_MTARGET_PRDATAS16;
input         M2_APB_MTARGET_PREADYS16;
input         M2_APB_MTARGET_PSLVERRS16;
input         M2_UART_CTS;
input         M2_UART_RXD;
input         MAC_1_MDI_F2M;
input         MMUART_2_RXD;
input         MMUART_3_RXD;
input         MMUART_4_RXD;
input  [58:3] MSS_INT_F2M;
input         PCIE_INT;
input         PHY_INTn;
input         PRESETN;
input         REFCLK;
input         REFCLK_N;
input         SD_DET;
input         SGMII_RX0_N;
input         SGMII_RX0_P;
input         SGMII_RX1_N;
input         SGMII_RX1_P;
input         SPI_0_DI;
input         SPI_1_DI;
input         UART0_RXD;
input         USB_CLK;
input         USB_DIR;
input         USB_NXT;
input         USB_OCn;
input         USER_BUTTON;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output        ADC_CSn;
output        ADC_SCK;
output [5:0]  CA;
output [31:0] CAPE_APB_MTARGET_PADDRS;
output        CAPE_APB_MTARGET_PENABLES;
output        CAPE_APB_MTARGET_PSELS1;
output [31:0] CAPE_APB_MTARGET_PWDATAS;
output        CAPE_APB_MTARGET_PWRITES;
output        CK;
output        CKE;
output        CK_N;
output        CS;
output        CSI_APB_MTARGET_PSELS2;
output [3:0]  DM;
output        EMMC_CLK;
output        EMMC_RSTN;
output [37:0] FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARADDR;
output [1:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARBURST;
output [3:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARCACHE;
output [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARID;
output [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARLEN;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARLOCK;
output [2:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARPROT;
output [3:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARQOS;
output [2:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARSIZE;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARVALID;
output [37:0] FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWADDR;
output [1:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWBURST;
output [3:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWCACHE;
output [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWID;
output [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWLEN;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWLOCK;
output [2:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWPROT;
output [3:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWQOS;
output [2:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWSIZE;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWVALID;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BREADY;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RREADY;
output [63:0] FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WDATA;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WLAST;
output [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WSTRB;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WVALID;
output        FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARREADY;
output        FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWREADY;
output [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BID;
output [1:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BRESP;
output        FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BVALID;
output [63:0] FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RDATA;
output [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RID;
output        FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RLAST;
output [1:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RRESP;
output        FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RVALID;
output        FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WREADY;
output [37:0] FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARADDR;
output [1:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARBURST;
output [3:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARCACHE;
output [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARID;
output [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARLEN;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARLOCK;
output [2:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARPROT;
output [3:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARQOS;
output [2:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARSIZE;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARVALID;
output [37:0] FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWADDR;
output [1:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWBURST;
output [3:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWCACHE;
output [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWID;
output [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWLEN;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWLOCK;
output [2:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWPROT;
output [3:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWQOS;
output [2:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWSIZE;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWVALID;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BREADY;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RREADY;
output [63:0] FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WDATA;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WLAST;
output [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WSTRB;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WVALID;
output        FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARREADY;
output        FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWREADY;
output [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BID;
output [1:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BRESP;
output        FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BVALID;
output [63:0] FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RDATA;
output [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RID;
output        FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RLAST;
output [1:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RRESP;
output        FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RVALID;
output        FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WREADY;
output        FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARREADY;
output        FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWREADY;
output [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BID;
output [1:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BRESP;
output        FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BVALID;
output [63:0] FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RDATA;
output [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RID;
output        FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RLAST;
output [1:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RRESP;
output        FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RVALID;
output        FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WREADY;
output [3:0]  FIC_3_APB_M_PSTRB;
output [27:0] GPIO_2_M2F;
output [27:0] GPIO_2_OE_M2F;
output        HSI_APB_MTARGET_PSELS4;
output        M2_APB_MTARGET_PSELS16;
output        M2_UART_RTS;
output        M2_UART_TXD;
output        M2_W_DISABLE1;
output        M2_W_DISABLE2;
output        MAC_1_MDC_M2F;
output        MAC_1_MDO_M2F;
output        MAC_1_MDO_OE_M2F;
output        MMUART_2_TXD;
output        MMUART_3_TXD;
output        MMUART_4_TXD;
output        MSS_DLL_LOCKS;
output        MSS_RESET_N_M2F;
output        ODT;
output        PHY_MDC;
output        RESET_N;
output        SD_CARD_CS;
output        SGMII_TX0_N;
output        SGMII_TX0_P;
output        SGMII_TX1_N;
output        SGMII_TX1_P;
output        SPI_0_CLK;
output        SPI_0_DO;
output        SPI_0_SS1;
output        SPI_1_CLK;
output        SPI_1_DO;
output        SPI_1_SS1;
output        UART0_TXD;
output        USB_STP;
output        VIO_ENABLE;
//--------------------------------------------------------------------
// Inout
//--------------------------------------------------------------------
inout         ADC_MISO;
inout         ADC_MOSI;
inout  [31:0] DQ;
inout  [3:0]  DQS;
inout  [3:0]  DQS_N;
inout         EMMC_CMD;
inout         EMMC_DATA0;
inout         EMMC_DATA1;
inout         EMMC_DATA2;
inout         EMMC_DATA3;
inout         EMMC_DATA4;
inout         EMMC_DATA5;
inout         EMMC_DATA6;
inout         EMMC_DATA7;
inout         I2C0_SCL;
inout         I2C0_SDA;
inout         I2C_1_SCL;
inout         I2C_1_SDA;
inout         PHY_MDIO;
inout         USB_DATA0;
inout         USB_DATA1;
inout         USB_DATA2;
inout         USB_DATA3;
inout         USB_DATA4;
inout         USB_DATA5;
inout         USB_DATA6;
inout         USB_DATA7;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire           ADC_CSn_net_0;
wire           ADC_IRQn;
wire           ADC_MISO;
wire           ADC_MOSI;
wire           ADC_SCK_net_0;
wire   [31:0]  APB_ARBITER_0_APB_MASTER_high_PADDR;
wire           APB_ARBITER_0_APB_MASTER_high_PENABLE;
wire   [31:0]  APB_ARBITER_0_APB_MASTER_high_PRDATA;
wire           APB_ARBITER_0_APB_MASTER_high_PREADY;
wire           APB_ARBITER_0_APB_MASTER_high_PSELx;
wire           APB_ARBITER_0_APB_MASTER_high_PSLVERR;
wire   [31:0]  APB_ARBITER_0_APB_MASTER_high_PWDATA;
wire           APB_ARBITER_0_APB_MASTER_high_PWRITE;
wire   [31:0]  APB_ARBITER_0_APB_MASTER_low_PADDR;
wire           APB_ARBITER_0_APB_MASTER_low_PENABLE;
wire   [31:0]  APB_ARBITER_0_APB_MASTER_low_PRDATA;
wire           APB_ARBITER_0_APB_MASTER_low_PREADY;
wire           APB_ARBITER_0_APB_MASTER_low_PSELx;
wire           APB_ARBITER_0_APB_MASTER_low_PSLVERR;
wire   [31:0]  APB_ARBITER_0_APB_MASTER_low_PWDATA;
wire           APB_ARBITER_0_APB_MASTER_low_PWRITE;
wire   [5:0]   CA_net_0;
wire   [31:0]  CAPE_APB_MTARGET_PADDR;
wire           CAPE_APB_MTARGET_PENABLE;
wire   [31:0]  CAPE_APB_MTARGET_PRDATAS1;
wire           CAPE_APB_MTARGET_PREADYS1;
wire           CAPE_APB_MTARGET_PSELx;
wire           CAPE_APB_MTARGET_PSLVERRS1;
wire   [31:0]  CAPE_APB_MTARGET_PWDATA;
wire           CAPE_APB_MTARGET_PWRITE;
wire           CK_net_0;
wire           CK_N_net_0;
wire           CKE_net_0;
wire           CS_net_0;
wire   [31:0]  CSI_APB_MTARGET_PRDATAS2;
wire           CSI_APB_MTARGET_PREADYS2;
wire           CSI_APB_MTARGET_PSELx;
wire           CSI_APB_MTARGET_PSLVERRS2;
wire   [3:0]   DM_net_0;
wire   [31:0]  DQ;
wire   [3:0]   DQS;
wire   [3:0]   DQS_N;
wire           EMMC_CLK_net_0;
wire           EMMC_CMD;
wire           EMMC_DATA0;
wire           EMMC_DATA1;
wire           EMMC_DATA2;
wire           EMMC_DATA3;
wire           EMMC_DATA4;
wire           EMMC_DATA5;
wire           EMMC_DATA6;
wire           EMMC_DATA7;
wire           EMMC_RSTN_net_0;
wire           EMMC_STRB;
wire           FIC_0_ACLK;
wire   [37:0]  FIC_0_AXI4_INITIATOR_ARADDR;
wire   [1:0]   FIC_0_AXI4_INITIATOR_ARBURST;
wire   [3:0]   FIC_0_AXI4_INITIATOR_ARCACHE;
wire   [7:0]   FIC_0_AXI4_INITIATOR_ARID;
wire   [7:0]   FIC_0_AXI4_INITIATOR_ARLEN;
wire           FIC_0_AXI4_INITIATOR_ARLOCK;
wire   [2:0]   FIC_0_AXI4_INITIATOR_ARPROT;
wire   [3:0]   FIC_0_AXI4_INITIATOR_ARQOS;
wire           FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARREADY;
wire   [2:0]   FIC_0_AXI4_INITIATOR_ARSIZE;
wire           FIC_0_AXI4_INITIATOR_ARVALID;
wire   [37:0]  FIC_0_AXI4_INITIATOR_AWADDR;
wire   [1:0]   FIC_0_AXI4_INITIATOR_AWBURST;
wire   [3:0]   FIC_0_AXI4_INITIATOR_AWCACHE;
wire   [7:0]   FIC_0_AXI4_INITIATOR_AWID;
wire   [7:0]   FIC_0_AXI4_INITIATOR_AWLEN;
wire           FIC_0_AXI4_INITIATOR_AWLOCK;
wire   [2:0]   FIC_0_AXI4_INITIATOR_AWPROT;
wire   [3:0]   FIC_0_AXI4_INITIATOR_AWQOS;
wire           FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWREADY;
wire   [2:0]   FIC_0_AXI4_INITIATOR_AWSIZE;
wire           FIC_0_AXI4_INITIATOR_AWVALID;
wire   [7:0]   FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BID;
wire           FIC_0_AXI4_INITIATOR_BREADY;
wire   [1:0]   FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BRESP;
wire           FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BVALID;
wire   [63:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RDATA;
wire   [7:0]   FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RID;
wire           FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RLAST;
wire           FIC_0_AXI4_INITIATOR_RREADY;
wire   [1:0]   FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RRESP;
wire           FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RVALID;
wire   [63:0]  FIC_0_AXI4_INITIATOR_WDATA;
wire           FIC_0_AXI4_INITIATOR_WLAST;
wire           FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WREADY;
wire   [7:0]   FIC_0_AXI4_INITIATOR_WSTRB;
wire           FIC_0_AXI4_INITIATOR_WVALID;
wire   [37:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARADDR;
wire   [1:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARBURST;
wire   [3:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARCACHE;
wire   [3:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARID;
wire   [7:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLEN;
wire           FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLOCK;
wire   [2:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARPROT;
wire   [3:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARQOS;
wire           FIC_0_AXI4_TARGET_ARREADY;
wire   [2:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARSIZE;
wire           FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARVALID;
wire   [37:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWADDR;
wire   [1:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWBURST;
wire   [3:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWCACHE;
wire   [3:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWID;
wire   [7:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLEN;
wire           FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLOCK;
wire   [2:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWPROT;
wire   [3:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWQOS;
wire           FIC_0_AXI4_TARGET_AWREADY;
wire   [2:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWSIZE;
wire           FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWVALID;
wire   [3:0]   FIC_0_AXI4_TARGET_BID;
wire           FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BREADY;
wire   [1:0]   FIC_0_AXI4_TARGET_BRESP;
wire           FIC_0_AXI4_TARGET_BVALID;
wire   [63:0]  FIC_0_AXI4_TARGET_RDATA;
wire   [3:0]   FIC_0_AXI4_TARGET_RID;
wire           FIC_0_AXI4_TARGET_RLAST;
wire           FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RREADY;
wire   [1:0]   FIC_0_AXI4_TARGET_RRESP;
wire           FIC_0_AXI4_TARGET_RVALID;
wire   [63:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WDATA;
wire           FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WLAST;
wire           FIC_0_AXI4_TARGET_WREADY;
wire   [7:0]   FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WSTRB;
wire           FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WVALID;
wire           FIC_1_ACLK;
wire   [37:0]  FIC_1_AXI4_INITIATOR_ARADDR;
wire   [1:0]   FIC_1_AXI4_INITIATOR_ARBURST;
wire   [3:0]   FIC_1_AXI4_INITIATOR_ARCACHE;
wire   [7:0]   FIC_1_AXI4_INITIATOR_ARID;
wire   [7:0]   FIC_1_AXI4_INITIATOR_ARLEN;
wire           FIC_1_AXI4_INITIATOR_ARLOCK;
wire   [2:0]   FIC_1_AXI4_INITIATOR_ARPROT;
wire   [3:0]   FIC_1_AXI4_INITIATOR_ARQOS;
wire           FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARREADY;
wire   [2:0]   FIC_1_AXI4_INITIATOR_ARSIZE;
wire           FIC_1_AXI4_INITIATOR_ARVALID;
wire   [37:0]  FIC_1_AXI4_INITIATOR_AWADDR;
wire   [1:0]   FIC_1_AXI4_INITIATOR_AWBURST;
wire   [3:0]   FIC_1_AXI4_INITIATOR_AWCACHE;
wire   [7:0]   FIC_1_AXI4_INITIATOR_AWID;
wire   [7:0]   FIC_1_AXI4_INITIATOR_AWLEN;
wire           FIC_1_AXI4_INITIATOR_AWLOCK;
wire   [2:0]   FIC_1_AXI4_INITIATOR_AWPROT;
wire   [3:0]   FIC_1_AXI4_INITIATOR_AWQOS;
wire           FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWREADY;
wire   [2:0]   FIC_1_AXI4_INITIATOR_AWSIZE;
wire           FIC_1_AXI4_INITIATOR_AWVALID;
wire   [7:0]   FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BID;
wire           FIC_1_AXI4_INITIATOR_BREADY;
wire   [1:0]   FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BRESP;
wire           FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BVALID;
wire   [63:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RDATA;
wire   [7:0]   FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RID;
wire           FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RLAST;
wire           FIC_1_AXI4_INITIATOR_RREADY;
wire   [1:0]   FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RRESP;
wire           FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RVALID;
wire   [63:0]  FIC_1_AXI4_INITIATOR_WDATA;
wire           FIC_1_AXI4_INITIATOR_WLAST;
wire           FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WREADY;
wire   [7:0]   FIC_1_AXI4_INITIATOR_WSTRB;
wire           FIC_1_AXI4_INITIATOR_WVALID;
wire   [37:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARADDR;
wire   [1:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARBURST;
wire   [3:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARCACHE;
wire   [3:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARID;
wire   [7:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLEN;
wire           FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLOCK;
wire   [2:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARPROT;
wire   [3:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARQOS;
wire           FIC_1_AXI4_TARGET_ARREADY;
wire   [2:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARSIZE;
wire           FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARVALID;
wire   [37:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWADDR;
wire   [1:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWBURST;
wire   [3:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWCACHE;
wire   [3:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWID;
wire   [7:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLEN;
wire           FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLOCK;
wire   [2:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWPROT;
wire   [3:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWQOS;
wire           FIC_1_AXI4_TARGET_AWREADY;
wire   [2:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWSIZE;
wire           FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWVALID;
wire   [3:0]   FIC_1_AXI4_TARGET_BID;
wire           FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BREADY;
wire   [1:0]   FIC_1_AXI4_TARGET_BRESP;
wire           FIC_1_AXI4_TARGET_BVALID;
wire   [63:0]  FIC_1_AXI4_TARGET_RDATA;
wire   [3:0]   FIC_1_AXI4_TARGET_RID;
wire           FIC_1_AXI4_TARGET_RLAST;
wire           FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RREADY;
wire   [1:0]   FIC_1_AXI4_TARGET_RRESP;
wire           FIC_1_AXI4_TARGET_RVALID;
wire   [63:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WDATA;
wire           FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WLAST;
wire           FIC_1_AXI4_TARGET_WREADY;
wire   [7:0]   FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WSTRB;
wire           FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WVALID;
wire           FIC_2_ACLK;
wire   [37:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARADDR;
wire   [1:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARBURST;
wire   [3:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARCACHE;
wire   [3:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARID;
wire   [7:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLEN;
wire           FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLOCK;
wire   [2:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARPROT;
wire   [3:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARQOS;
wire           FIC_2_AXI4_TARGET_ARREADY;
wire   [2:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARSIZE;
wire           FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARVALID;
wire   [37:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWADDR;
wire   [1:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWBURST;
wire   [3:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWCACHE;
wire   [3:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWID;
wire   [7:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLEN;
wire           FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLOCK;
wire   [2:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWPROT;
wire   [3:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWQOS;
wire           FIC_2_AXI4_TARGET_AWREADY;
wire   [2:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWSIZE;
wire           FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWVALID;
wire   [3:0]   FIC_2_AXI4_TARGET_BID;
wire           FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BREADY;
wire   [1:0]   FIC_2_AXI4_TARGET_BRESP;
wire           FIC_2_AXI4_TARGET_BVALID;
wire   [63:0]  FIC_2_AXI4_TARGET_RDATA;
wire   [3:0]   FIC_2_AXI4_TARGET_RID;
wire           FIC_2_AXI4_TARGET_RLAST;
wire           FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RREADY;
wire   [1:0]   FIC_2_AXI4_TARGET_RRESP;
wire           FIC_2_AXI4_TARGET_RVALID;
wire   [63:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WDATA;
wire           FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WLAST;
wire           FIC_2_AXI4_TARGET_WREADY;
wire   [7:0]   FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WSTRB;
wire           FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WVALID;
wire   [3:0]   FIC_3_APB_M_PSTRB_net_0;
wire           FIC_3_PCLK;
wire   [27:27] GPIO_2_F2M_slice_0;
wire   [26:26] GPIO_2_F2M_slice_1;
wire   [25:25] GPIO_2_F2M_slice_2;
wire   [24:24] GPIO_2_F2M_slice_3;
wire   [23:23] GPIO_2_F2M_slice_4;
wire   [22:22] GPIO_2_F2M_slice_5;
wire   [21:21] GPIO_2_F2M_slice_6;
wire   [20:20] GPIO_2_F2M_slice_7;
wire   [19:19] GPIO_2_F2M_slice_8;
wire   [18:18] GPIO_2_F2M_slice_9;
wire   [17:17] GPIO_2_F2M_slice_10;
wire   [16:16] GPIO_2_F2M_slice_11;
wire   [15:15] GPIO_2_F2M_slice_12;
wire   [14:14] GPIO_2_F2M_slice_13;
wire   [13:13] GPIO_2_F2M_slice_14;
wire   [12:12] GPIO_2_F2M_slice_15;
wire   [11:11] GPIO_2_F2M_slice_16;
wire   [10:10] GPIO_2_F2M_slice_17;
wire   [9:9]   GPIO_2_F2M_slice_18;
wire   [8:8]   GPIO_2_F2M_slice_19;
wire   [7:7]   GPIO_2_F2M_slice_20;
wire   [6:6]   GPIO_2_F2M_slice_21;
wire   [5:5]   GPIO_2_F2M_slice_22;
wire   [4:4]   GPIO_2_F2M_slice_23;
wire   [3:3]   GPIO_2_F2M_slice_24;
wire   [2:2]   GPIO_2_F2M_slice_25;
wire   [1:1]   GPIO_2_F2M_slice_26;
wire   [0:0]   GPIO_2_F2M_slice_27;
wire           GPIO_2_M2F_net_0;
wire           GPIO_2_M2F_0;
wire           GPIO_2_M2F_1;
wire           GPIO_2_M2F_2;
wire           GPIO_2_M2F_3;
wire           GPIO_2_M2F_4;
wire           GPIO_2_M2F_5;
wire           GPIO_2_M2F_6;
wire           GPIO_2_M2F_7;
wire           GPIO_2_M2F_8;
wire           GPIO_2_M2F_9;
wire           GPIO_2_M2F_10;
wire           GPIO_2_M2F_11;
wire           GPIO_2_M2F_12;
wire           GPIO_2_M2F_13;
wire           GPIO_2_M2F_14;
wire           GPIO_2_M2F_15;
wire           GPIO_2_M2F_16;
wire           GPIO_2_M2F_17;
wire           GPIO_2_M2F_18;
wire           GPIO_2_M2F_19;
wire           GPIO_2_M2F_20;
wire           GPIO_2_M2F_21;
wire           GPIO_2_M2F_22;
wire           GPIO_2_M2F_23;
wire           GPIO_2_M2F_24;
wire           GPIO_2_M2F_25;
wire           GPIO_2_M2F_26;
wire           GPIO_2_OE_M2F_net_0;
wire           GPIO_2_OE_M2F_0;
wire           GPIO_2_OE_M2F_1;
wire           GPIO_2_OE_M2F_2;
wire           GPIO_2_OE_M2F_3;
wire           GPIO_2_OE_M2F_4;
wire           GPIO_2_OE_M2F_5;
wire           GPIO_2_OE_M2F_6;
wire           GPIO_2_OE_M2F_7;
wire           GPIO_2_OE_M2F_8;
wire           GPIO_2_OE_M2F_9;
wire           GPIO_2_OE_M2F_10;
wire           GPIO_2_OE_M2F_11;
wire           GPIO_2_OE_M2F_12;
wire           GPIO_2_OE_M2F_13;
wire           GPIO_2_OE_M2F_14;
wire           GPIO_2_OE_M2F_15;
wire           GPIO_2_OE_M2F_16;
wire           GPIO_2_OE_M2F_17;
wire           GPIO_2_OE_M2F_18;
wire           GPIO_2_OE_M2F_19;
wire           GPIO_2_OE_M2F_20;
wire           GPIO_2_OE_M2F_21;
wire           GPIO_2_OE_M2F_22;
wire           GPIO_2_OE_M2F_23;
wire           GPIO_2_OE_M2F_24;
wire           GPIO_2_OE_M2F_25;
wire           GPIO_2_OE_M2F_26;
wire   [31:0]  HSI_APB_MTARGET_PRDATAS4;
wire           HSI_APB_MTARGET_PREADYS4;
wire           HSI_APB_MTARGET_PSELx;
wire           HSI_APB_MTARGET_PSLVERRS4;
wire           I2C0_SCL;
wire           I2C0_SCL_BIBUF_Y;
wire           I2C0_SDA;
wire           I2C0_SDA_BIBUF_Y;
wire           I2C_1_SCL;
wire           I2C_1_SDA;
wire           IHC_SUBSYSTEM_0_E51_IRQ;
wire           IHC_SUBSYSTEM_0_U54_1_IRQ;
wire           IHC_SUBSYSTEM_0_U54_2_IRQ;
wire           IHC_SUBSYSTEM_0_U54_3_IRQ;
wire           IHC_SUBSYSTEM_0_U54_4_IRQ;
wire   [31:0]  M2_APB_MTARGET_PRDATAS16;
wire           M2_APB_MTARGET_PREADYS16;
wire           M2_APB_MTARGET_PSELx;
wire           M2_APB_MTARGET_PSLVERRS16;
wire           M2_UART_CTS;
wire           M2_UART_RTS_net_0;
wire           M2_UART_RXD;
wire           M2_UART_TXD_net_0;
wire           M2_W_DISABLE1_net_0;
wire           M2_W_DISABLE2_net_0;
wire           MAC_1_MDC_M2F_net_0;
wire           MAC_1_MDI_F2M;
wire           MAC_1_MDO_M2F_net_0;
wire           MAC_1_MDO_OE_M2F_net_0;
wire           MMUART_2_RXD;
wire           MMUART_2_TXD_net_0;
wire           MMUART_3_RXD;
wire           MMUART_3_TXD_net_0;
wire           MMUART_4_RXD;
wire           MMUART_4_TXD_net_0;
wire           MSS_DLL_LOCKS_net_0;
wire   [58:3]  MSS_INT_F2M;
wire           MSS_RESET_N_M2F_net_0;
wire           ODT_net_0;
wire           PCIE_INT;
wire           PF_SOC_MSS_FIC_0_DLL_LOCK_M2F;
wire           PF_SOC_MSS_FIC_1_DLL_LOCK_M2F;
wire           PF_SOC_MSS_FIC_2_DLL_LOCK_M2F;
wire   [31:0]  PF_SOC_MSS_FIC_3_APB_INITIATOR_PADDR;
wire           PF_SOC_MSS_FIC_3_APB_INITIATOR_PENABLE;
wire   [31:0]  PF_SOC_MSS_FIC_3_APB_INITIATOR_PRDATA;
wire           PF_SOC_MSS_FIC_3_APB_INITIATOR_PREADY;
wire           PF_SOC_MSS_FIC_3_APB_INITIATOR_PSELx;
wire           PF_SOC_MSS_FIC_3_APB_INITIATOR_PSLVERR;
wire   [31:0]  PF_SOC_MSS_FIC_3_APB_INITIATOR_PWDATA;
wire           PF_SOC_MSS_FIC_3_APB_INITIATOR_PWRITE;
wire           PF_SOC_MSS_FIC_3_DLL_LOCK_M2F;
wire           PF_SOC_MSS_I2C_0_SCL_OE_M2F;
wire           PF_SOC_MSS_I2C_0_SDA_OE_M2F;
wire           PHY_INTn;
wire           PHY_MDC_net_0;
wire           PHY_MDIO;
wire           PRESETN;
wire           REFCLK;
wire           REFCLK_N;
wire           RESET_N_net_0;
wire           SD_CARD_CS_net_0;
wire           SD_DET;
wire           SGMII_RX0_N;
wire           SGMII_RX0_P;
wire           SGMII_RX1_N;
wire           SGMII_RX1_P;
wire           SGMII_TX0_N_net_0;
wire           SGMII_TX0_P_net_0;
wire           SGMII_TX1_N_net_0;
wire           SGMII_TX1_P_net_0;
wire           SPI_0_CLK_net_0;
wire           SPI_0_DI;
wire           SPI_0_DO_net_0;
wire           SPI_0_SS1_net_0;
wire           SPI_1_CLK_net_0;
wire           SPI_1_DI;
wire           SPI_1_DO_net_0;
wire           SPI_1_SS1_net_0;
wire           UART0_RXD;
wire           UART0_TXD_net_0;
wire           USB_CLK;
wire           USB_DATA0;
wire           USB_DATA1;
wire           USB_DATA2;
wire           USB_DATA3;
wire           USB_DATA4;
wire           USB_DATA5;
wire           USB_DATA6;
wire           USB_DATA7;
wire           USB_DIR;
wire           USB_NXT;
wire           USB_OCn;
wire           USB_STP_net_0;
wire           USER_BUTTON;
wire           VIO_ENABLE_net_0;
wire           USB_STP_net_1;
wire           UART0_TXD_net_1;
wire           M2_UART_TXD_net_1;
wire           M2_UART_RTS_net_1;
wire           MSS_DLL_LOCKS_net_1;
wire           RESET_N_net_1;
wire           ODT_net_1;
wire           CKE_net_1;
wire           CS_net_1;
wire           CK_net_1;
wire           CK_N_net_1;
wire           SGMII_TX0_P_net_1;
wire           SGMII_TX0_N_net_1;
wire           SGMII_TX1_P_net_1;
wire           SGMII_TX1_N_net_1;
wire   [5:0]   CA_net_1;
wire   [3:0]   DM_net_1;
wire           SD_CARD_CS_net_1;
wire   [0:0]   GPIO_2_M2F_26_net_0;
wire   [10:10] GPIO_2_M2F_16_net_0;
wire   [11:11] GPIO_2_M2F_15_net_0;
wire   [12:12] GPIO_2_M2F_14_net_0;
wire   [13:13] GPIO_2_M2F_13_net_0;
wire   [14:14] GPIO_2_M2F_12_net_0;
wire   [15:15] GPIO_2_M2F_11_net_0;
wire   [16:16] GPIO_2_M2F_10_net_0;
wire   [17:17] GPIO_2_M2F_9_net_0;
wire   [18:18] GPIO_2_M2F_8_net_0;
wire   [19:19] GPIO_2_M2F_7_net_0;
wire   [1:1]   GPIO_2_M2F_25_net_0;
wire   [20:20] GPIO_2_M2F_6_net_0;
wire   [21:21] GPIO_2_M2F_5_net_0;
wire   [22:22] GPIO_2_M2F_4_net_0;
wire   [23:23] GPIO_2_M2F_3_net_0;
wire   [24:24] GPIO_2_M2F_2_net_0;
wire   [25:25] GPIO_2_M2F_1_net_0;
wire   [26:26] GPIO_2_M2F_0_net_0;
wire   [27:27] GPIO_2_M2F_net_1;
wire   [2:2]   GPIO_2_M2F_24_net_0;
wire   [3:3]   GPIO_2_M2F_23_net_0;
wire   [4:4]   GPIO_2_M2F_22_net_0;
wire   [5:5]   GPIO_2_M2F_21_net_0;
wire   [6:6]   GPIO_2_M2F_20_net_0;
wire   [7:7]   GPIO_2_M2F_19_net_0;
wire   [8:8]   GPIO_2_M2F_18_net_0;
wire   [9:9]   GPIO_2_M2F_17_net_0;
wire   [0:0]   GPIO_2_OE_M2F_26_net_0;
wire   [10:10] GPIO_2_OE_M2F_16_net_0;
wire   [11:11] GPIO_2_OE_M2F_15_net_0;
wire   [12:12] GPIO_2_OE_M2F_14_net_0;
wire   [13:13] GPIO_2_OE_M2F_13_net_0;
wire   [14:14] GPIO_2_OE_M2F_12_net_0;
wire   [15:15] GPIO_2_OE_M2F_11_net_0;
wire   [16:16] GPIO_2_OE_M2F_10_net_0;
wire   [17:17] GPIO_2_OE_M2F_9_net_0;
wire   [18:18] GPIO_2_OE_M2F_8_net_0;
wire   [19:19] GPIO_2_OE_M2F_7_net_0;
wire   [1:1]   GPIO_2_OE_M2F_25_net_0;
wire   [20:20] GPIO_2_OE_M2F_6_net_0;
wire   [21:21] GPIO_2_OE_M2F_5_net_0;
wire   [22:22] GPIO_2_OE_M2F_4_net_0;
wire   [23:23] GPIO_2_OE_M2F_3_net_0;
wire   [24:24] GPIO_2_OE_M2F_2_net_0;
wire   [25:25] GPIO_2_OE_M2F_1_net_0;
wire   [26:26] GPIO_2_OE_M2F_0_net_0;
wire   [27:27] GPIO_2_OE_M2F_net_1;
wire   [2:2]   GPIO_2_OE_M2F_24_net_0;
wire   [3:3]   GPIO_2_OE_M2F_23_net_0;
wire   [4:4]   GPIO_2_OE_M2F_22_net_0;
wire   [5:5]   GPIO_2_OE_M2F_21_net_0;
wire   [6:6]   GPIO_2_OE_M2F_20_net_0;
wire   [7:7]   GPIO_2_OE_M2F_19_net_0;
wire   [8:8]   GPIO_2_OE_M2F_18_net_0;
wire   [9:9]   GPIO_2_OE_M2F_17_net_0;
wire           ADC_CSn_net_1;
wire           ADC_SCK_net_1;
wire           MMUART_2_TXD_net_1;
wire           MMUART_3_TXD_net_1;
wire           MMUART_4_TXD_net_1;
wire           PHY_MDC_net_1;
wire           M2_W_DISABLE1_net_1;
wire           M2_W_DISABLE2_net_1;
wire           MAC_1_MDO_OE_M2F_net_1;
wire           MAC_1_MDC_M2F_net_1;
wire           MAC_1_MDO_M2F_net_1;
wire           EMMC_CLK_net_1;
wire           EMMC_RSTN_net_1;
wire           VIO_ENABLE_net_1;
wire           FIC_2_AXI4_TARGET_AWREADY_net_0;
wire           FIC_2_AXI4_TARGET_WREADY_net_0;
wire   [3:0]   FIC_2_AXI4_TARGET_BID_net_0;
wire   [1:0]   FIC_2_AXI4_TARGET_BRESP_net_0;
wire           FIC_2_AXI4_TARGET_BVALID_net_0;
wire           FIC_2_AXI4_TARGET_ARREADY_net_0;
wire   [3:0]   FIC_2_AXI4_TARGET_RID_net_0;
wire   [63:0]  FIC_2_AXI4_TARGET_RDATA_net_0;
wire   [1:0]   FIC_2_AXI4_TARGET_RRESP_net_0;
wire           FIC_2_AXI4_TARGET_RLAST_net_0;
wire           FIC_2_AXI4_TARGET_RVALID_net_0;
wire           FIC_1_AXI4_TARGET_AWREADY_net_0;
wire           FIC_1_AXI4_TARGET_WREADY_net_0;
wire   [3:0]   FIC_1_AXI4_TARGET_BID_net_0;
wire   [1:0]   FIC_1_AXI4_TARGET_BRESP_net_0;
wire           FIC_1_AXI4_TARGET_BVALID_net_0;
wire           FIC_1_AXI4_TARGET_ARREADY_net_0;
wire   [3:0]   FIC_1_AXI4_TARGET_RID_net_0;
wire   [63:0]  FIC_1_AXI4_TARGET_RDATA_net_0;
wire   [1:0]   FIC_1_AXI4_TARGET_RRESP_net_0;
wire           FIC_1_AXI4_TARGET_RLAST_net_0;
wire           FIC_1_AXI4_TARGET_RVALID_net_0;
wire           FIC_0_AXI4_TARGET_AWREADY_net_0;
wire           FIC_0_AXI4_TARGET_WREADY_net_0;
wire   [3:0]   FIC_0_AXI4_TARGET_BID_net_0;
wire   [1:0]   FIC_0_AXI4_TARGET_BRESP_net_0;
wire           FIC_0_AXI4_TARGET_BVALID_net_0;
wire           FIC_0_AXI4_TARGET_ARREADY_net_0;
wire   [3:0]   FIC_0_AXI4_TARGET_RID_net_0;
wire   [63:0]  FIC_0_AXI4_TARGET_RDATA_net_0;
wire   [1:0]   FIC_0_AXI4_TARGET_RRESP_net_0;
wire           FIC_0_AXI4_TARGET_RLAST_net_0;
wire           FIC_0_AXI4_TARGET_RVALID_net_0;
wire   [31:0]  CAPE_APB_MTARGET_PADDR_net_0;
wire           CAPE_APB_MTARGET_PSELx_net_0;
wire           CAPE_APB_MTARGET_PENABLE_net_0;
wire           CAPE_APB_MTARGET_PWRITE_net_0;
wire   [31:0]  CAPE_APB_MTARGET_PWDATA_net_0;
wire           CSI_APB_MTARGET_PSELx_net_0;
wire           HSI_APB_MTARGET_PSELx_net_0;
wire           M2_APB_MTARGET_PSELx_net_0;
wire           MSS_RESET_N_M2F_net_1;
wire   [3:0]   FIC_3_APB_M_PSTRB_net_1;
wire   [7:0]   FIC_0_AXI4_INITIATOR_AWID_net_0;
wire   [37:0]  FIC_0_AXI4_INITIATOR_AWADDR_net_0;
wire   [7:0]   FIC_0_AXI4_INITIATOR_AWLEN_net_0;
wire   [2:0]   FIC_0_AXI4_INITIATOR_AWSIZE_net_0;
wire   [1:0]   FIC_0_AXI4_INITIATOR_AWBURST_net_0;
wire           FIC_0_AXI4_INITIATOR_AWLOCK_net_0;
wire   [3:0]   FIC_0_AXI4_INITIATOR_AWQOS_net_0;
wire   [3:0]   FIC_0_AXI4_INITIATOR_AWCACHE_net_0;
wire   [2:0]   FIC_0_AXI4_INITIATOR_AWPROT_net_0;
wire           FIC_0_AXI4_INITIATOR_AWVALID_net_0;
wire   [63:0]  FIC_0_AXI4_INITIATOR_WDATA_net_0;
wire   [7:0]   FIC_0_AXI4_INITIATOR_WSTRB_net_0;
wire           FIC_0_AXI4_INITIATOR_WLAST_net_0;
wire           FIC_0_AXI4_INITIATOR_WVALID_net_0;
wire           FIC_0_AXI4_INITIATOR_BREADY_net_0;
wire   [7:0]   FIC_0_AXI4_INITIATOR_ARID_net_0;
wire   [37:0]  FIC_0_AXI4_INITIATOR_ARADDR_net_0;
wire   [7:0]   FIC_0_AXI4_INITIATOR_ARLEN_net_0;
wire   [2:0]   FIC_0_AXI4_INITIATOR_ARSIZE_net_0;
wire   [1:0]   FIC_0_AXI4_INITIATOR_ARBURST_net_0;
wire           FIC_0_AXI4_INITIATOR_ARLOCK_net_0;
wire   [3:0]   FIC_0_AXI4_INITIATOR_ARQOS_net_0;
wire   [3:0]   FIC_0_AXI4_INITIATOR_ARCACHE_net_0;
wire   [2:0]   FIC_0_AXI4_INITIATOR_ARPROT_net_0;
wire           FIC_0_AXI4_INITIATOR_ARVALID_net_0;
wire           FIC_0_AXI4_INITIATOR_RREADY_net_0;
wire   [7:0]   FIC_1_AXI4_INITIATOR_AWID_net_0;
wire   [37:0]  FIC_1_AXI4_INITIATOR_AWADDR_net_0;
wire   [7:0]   FIC_1_AXI4_INITIATOR_AWLEN_net_0;
wire   [2:0]   FIC_1_AXI4_INITIATOR_AWSIZE_net_0;
wire   [1:0]   FIC_1_AXI4_INITIATOR_AWBURST_net_0;
wire           FIC_1_AXI4_INITIATOR_AWLOCK_net_0;
wire   [3:0]   FIC_1_AXI4_INITIATOR_AWQOS_net_0;
wire   [3:0]   FIC_1_AXI4_INITIATOR_AWCACHE_net_0;
wire   [2:0]   FIC_1_AXI4_INITIATOR_AWPROT_net_0;
wire           FIC_1_AXI4_INITIATOR_AWVALID_net_0;
wire   [63:0]  FIC_1_AXI4_INITIATOR_WDATA_net_0;
wire   [7:0]   FIC_1_AXI4_INITIATOR_WSTRB_net_0;
wire           FIC_1_AXI4_INITIATOR_WLAST_net_0;
wire           FIC_1_AXI4_INITIATOR_WVALID_net_0;
wire           FIC_1_AXI4_INITIATOR_BREADY_net_0;
wire   [7:0]   FIC_1_AXI4_INITIATOR_ARID_net_0;
wire   [37:0]  FIC_1_AXI4_INITIATOR_ARADDR_net_0;
wire   [7:0]   FIC_1_AXI4_INITIATOR_ARLEN_net_0;
wire   [2:0]   FIC_1_AXI4_INITIATOR_ARSIZE_net_0;
wire   [1:0]   FIC_1_AXI4_INITIATOR_ARBURST_net_0;
wire           FIC_1_AXI4_INITIATOR_ARLOCK_net_0;
wire   [3:0]   FIC_1_AXI4_INITIATOR_ARQOS_net_0;
wire   [3:0]   FIC_1_AXI4_INITIATOR_ARCACHE_net_0;
wire   [2:0]   FIC_1_AXI4_INITIATOR_ARPROT_net_0;
wire           FIC_1_AXI4_INITIATOR_ARVALID_net_0;
wire           FIC_1_AXI4_INITIATOR_RREADY_net_0;
wire           SPI_0_CLK_net_1;
wire           SPI_0_DO_net_1;
wire           SPI_0_SS1_net_1;
wire           SPI_1_SS1_net_1;
wire           SPI_1_CLK_net_1;
wire           SPI_1_DO_net_1;
wire   [27:0]  GPIO_2_F2M;
wire   [63:0]  MSS_INT_F2M_net_0;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire           GND_net;
wire           VCC_net;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net    = 1'b0;
assign VCC_net    = 1'b1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign USB_STP_net_1                                  = USB_STP_net_0;
assign USB_STP                                        = USB_STP_net_1;
assign UART0_TXD_net_1                                = UART0_TXD_net_0;
assign UART0_TXD                                      = UART0_TXD_net_1;
assign M2_UART_TXD_net_1                              = M2_UART_TXD_net_0;
assign M2_UART_TXD                                    = M2_UART_TXD_net_1;
assign M2_UART_RTS_net_1                              = M2_UART_RTS_net_0;
assign M2_UART_RTS                                    = M2_UART_RTS_net_1;
assign MSS_DLL_LOCKS_net_1                            = MSS_DLL_LOCKS_net_0;
assign MSS_DLL_LOCKS                                  = MSS_DLL_LOCKS_net_1;
assign RESET_N_net_1                                  = RESET_N_net_0;
assign RESET_N                                        = RESET_N_net_1;
assign ODT_net_1                                      = ODT_net_0;
assign ODT                                            = ODT_net_1;
assign CKE_net_1                                      = CKE_net_0;
assign CKE                                            = CKE_net_1;
assign CS_net_1                                       = CS_net_0;
assign CS                                             = CS_net_1;
assign CK_net_1                                       = CK_net_0;
assign CK                                             = CK_net_1;
assign CK_N_net_1                                     = CK_N_net_0;
assign CK_N                                           = CK_N_net_1;
assign SGMII_TX0_P_net_1                              = SGMII_TX0_P_net_0;
assign SGMII_TX0_P                                    = SGMII_TX0_P_net_1;
assign SGMII_TX0_N_net_1                              = SGMII_TX0_N_net_0;
assign SGMII_TX0_N                                    = SGMII_TX0_N_net_1;
assign SGMII_TX1_P_net_1                              = SGMII_TX1_P_net_0;
assign SGMII_TX1_P                                    = SGMII_TX1_P_net_1;
assign SGMII_TX1_N_net_1                              = SGMII_TX1_N_net_0;
assign SGMII_TX1_N                                    = SGMII_TX1_N_net_1;
assign CA_net_1                                       = CA_net_0;
assign CA[5:0]                                        = CA_net_1;
assign DM_net_1                                       = DM_net_0;
assign DM[3:0]                                        = DM_net_1;
assign SD_CARD_CS_net_1                               = SD_CARD_CS_net_0;
assign SD_CARD_CS                                     = SD_CARD_CS_net_1;
assign GPIO_2_M2F_26_net_0[0]                         = GPIO_2_M2F_26;
assign GPIO_2_M2F[0:0]                                = GPIO_2_M2F_26_net_0[0];
assign GPIO_2_M2F_16_net_0[10]                        = GPIO_2_M2F_16;
assign GPIO_2_M2F[10:10]                              = GPIO_2_M2F_16_net_0[10];
assign GPIO_2_M2F_15_net_0[11]                        = GPIO_2_M2F_15;
assign GPIO_2_M2F[11:11]                              = GPIO_2_M2F_15_net_0[11];
assign GPIO_2_M2F_14_net_0[12]                        = GPIO_2_M2F_14;
assign GPIO_2_M2F[12:12]                              = GPIO_2_M2F_14_net_0[12];
assign GPIO_2_M2F_13_net_0[13]                        = GPIO_2_M2F_13;
assign GPIO_2_M2F[13:13]                              = GPIO_2_M2F_13_net_0[13];
assign GPIO_2_M2F_12_net_0[14]                        = GPIO_2_M2F_12;
assign GPIO_2_M2F[14:14]                              = GPIO_2_M2F_12_net_0[14];
assign GPIO_2_M2F_11_net_0[15]                        = GPIO_2_M2F_11;
assign GPIO_2_M2F[15:15]                              = GPIO_2_M2F_11_net_0[15];
assign GPIO_2_M2F_10_net_0[16]                        = GPIO_2_M2F_10;
assign GPIO_2_M2F[16:16]                              = GPIO_2_M2F_10_net_0[16];
assign GPIO_2_M2F_9_net_0[17]                         = GPIO_2_M2F_9;
assign GPIO_2_M2F[17:17]                              = GPIO_2_M2F_9_net_0[17];
assign GPIO_2_M2F_8_net_0[18]                         = GPIO_2_M2F_8;
assign GPIO_2_M2F[18:18]                              = GPIO_2_M2F_8_net_0[18];
assign GPIO_2_M2F_7_net_0[19]                         = GPIO_2_M2F_7;
assign GPIO_2_M2F[19:19]                              = GPIO_2_M2F_7_net_0[19];
assign GPIO_2_M2F_25_net_0[1]                         = GPIO_2_M2F_25;
assign GPIO_2_M2F[1:1]                                = GPIO_2_M2F_25_net_0[1];
assign GPIO_2_M2F_6_net_0[20]                         = GPIO_2_M2F_6;
assign GPIO_2_M2F[20:20]                              = GPIO_2_M2F_6_net_0[20];
assign GPIO_2_M2F_5_net_0[21]                         = GPIO_2_M2F_5;
assign GPIO_2_M2F[21:21]                              = GPIO_2_M2F_5_net_0[21];
assign GPIO_2_M2F_4_net_0[22]                         = GPIO_2_M2F_4;
assign GPIO_2_M2F[22:22]                              = GPIO_2_M2F_4_net_0[22];
assign GPIO_2_M2F_3_net_0[23]                         = GPIO_2_M2F_3;
assign GPIO_2_M2F[23:23]                              = GPIO_2_M2F_3_net_0[23];
assign GPIO_2_M2F_2_net_0[24]                         = GPIO_2_M2F_2;
assign GPIO_2_M2F[24:24]                              = GPIO_2_M2F_2_net_0[24];
assign GPIO_2_M2F_1_net_0[25]                         = GPIO_2_M2F_1;
assign GPIO_2_M2F[25:25]                              = GPIO_2_M2F_1_net_0[25];
assign GPIO_2_M2F_0_net_0[26]                         = GPIO_2_M2F_0;
assign GPIO_2_M2F[26:26]                              = GPIO_2_M2F_0_net_0[26];
assign GPIO_2_M2F_net_1[27]                           = GPIO_2_M2F_net_0;
assign GPIO_2_M2F[27:27]                              = GPIO_2_M2F_net_1[27];
assign GPIO_2_M2F_24_net_0[2]                         = GPIO_2_M2F_24;
assign GPIO_2_M2F[2:2]                                = GPIO_2_M2F_24_net_0[2];
assign GPIO_2_M2F_23_net_0[3]                         = GPIO_2_M2F_23;
assign GPIO_2_M2F[3:3]                                = GPIO_2_M2F_23_net_0[3];
assign GPIO_2_M2F_22_net_0[4]                         = GPIO_2_M2F_22;
assign GPIO_2_M2F[4:4]                                = GPIO_2_M2F_22_net_0[4];
assign GPIO_2_M2F_21_net_0[5]                         = GPIO_2_M2F_21;
assign GPIO_2_M2F[5:5]                                = GPIO_2_M2F_21_net_0[5];
assign GPIO_2_M2F_20_net_0[6]                         = GPIO_2_M2F_20;
assign GPIO_2_M2F[6:6]                                = GPIO_2_M2F_20_net_0[6];
assign GPIO_2_M2F_19_net_0[7]                         = GPIO_2_M2F_19;
assign GPIO_2_M2F[7:7]                                = GPIO_2_M2F_19_net_0[7];
assign GPIO_2_M2F_18_net_0[8]                         = GPIO_2_M2F_18;
assign GPIO_2_M2F[8:8]                                = GPIO_2_M2F_18_net_0[8];
assign GPIO_2_M2F_17_net_0[9]                         = GPIO_2_M2F_17;
assign GPIO_2_M2F[9:9]                                = GPIO_2_M2F_17_net_0[9];
assign GPIO_2_OE_M2F_26_net_0[0]                      = GPIO_2_OE_M2F_26;
assign GPIO_2_OE_M2F[0:0]                             = GPIO_2_OE_M2F_26_net_0[0];
assign GPIO_2_OE_M2F_16_net_0[10]                     = GPIO_2_OE_M2F_16;
assign GPIO_2_OE_M2F[10:10]                           = GPIO_2_OE_M2F_16_net_0[10];
assign GPIO_2_OE_M2F_15_net_0[11]                     = GPIO_2_OE_M2F_15;
assign GPIO_2_OE_M2F[11:11]                           = GPIO_2_OE_M2F_15_net_0[11];
assign GPIO_2_OE_M2F_14_net_0[12]                     = GPIO_2_OE_M2F_14;
assign GPIO_2_OE_M2F[12:12]                           = GPIO_2_OE_M2F_14_net_0[12];
assign GPIO_2_OE_M2F_13_net_0[13]                     = GPIO_2_OE_M2F_13;
assign GPIO_2_OE_M2F[13:13]                           = GPIO_2_OE_M2F_13_net_0[13];
assign GPIO_2_OE_M2F_12_net_0[14]                     = GPIO_2_OE_M2F_12;
assign GPIO_2_OE_M2F[14:14]                           = GPIO_2_OE_M2F_12_net_0[14];
assign GPIO_2_OE_M2F_11_net_0[15]                     = GPIO_2_OE_M2F_11;
assign GPIO_2_OE_M2F[15:15]                           = GPIO_2_OE_M2F_11_net_0[15];
assign GPIO_2_OE_M2F_10_net_0[16]                     = GPIO_2_OE_M2F_10;
assign GPIO_2_OE_M2F[16:16]                           = GPIO_2_OE_M2F_10_net_0[16];
assign GPIO_2_OE_M2F_9_net_0[17]                      = GPIO_2_OE_M2F_9;
assign GPIO_2_OE_M2F[17:17]                           = GPIO_2_OE_M2F_9_net_0[17];
assign GPIO_2_OE_M2F_8_net_0[18]                      = GPIO_2_OE_M2F_8;
assign GPIO_2_OE_M2F[18:18]                           = GPIO_2_OE_M2F_8_net_0[18];
assign GPIO_2_OE_M2F_7_net_0[19]                      = GPIO_2_OE_M2F_7;
assign GPIO_2_OE_M2F[19:19]                           = GPIO_2_OE_M2F_7_net_0[19];
assign GPIO_2_OE_M2F_25_net_0[1]                      = GPIO_2_OE_M2F_25;
assign GPIO_2_OE_M2F[1:1]                             = GPIO_2_OE_M2F_25_net_0[1];
assign GPIO_2_OE_M2F_6_net_0[20]                      = GPIO_2_OE_M2F_6;
assign GPIO_2_OE_M2F[20:20]                           = GPIO_2_OE_M2F_6_net_0[20];
assign GPIO_2_OE_M2F_5_net_0[21]                      = GPIO_2_OE_M2F_5;
assign GPIO_2_OE_M2F[21:21]                           = GPIO_2_OE_M2F_5_net_0[21];
assign GPIO_2_OE_M2F_4_net_0[22]                      = GPIO_2_OE_M2F_4;
assign GPIO_2_OE_M2F[22:22]                           = GPIO_2_OE_M2F_4_net_0[22];
assign GPIO_2_OE_M2F_3_net_0[23]                      = GPIO_2_OE_M2F_3;
assign GPIO_2_OE_M2F[23:23]                           = GPIO_2_OE_M2F_3_net_0[23];
assign GPIO_2_OE_M2F_2_net_0[24]                      = GPIO_2_OE_M2F_2;
assign GPIO_2_OE_M2F[24:24]                           = GPIO_2_OE_M2F_2_net_0[24];
assign GPIO_2_OE_M2F_1_net_0[25]                      = GPIO_2_OE_M2F_1;
assign GPIO_2_OE_M2F[25:25]                           = GPIO_2_OE_M2F_1_net_0[25];
assign GPIO_2_OE_M2F_0_net_0[26]                      = GPIO_2_OE_M2F_0;
assign GPIO_2_OE_M2F[26:26]                           = GPIO_2_OE_M2F_0_net_0[26];
assign GPIO_2_OE_M2F_net_1[27]                        = GPIO_2_OE_M2F_net_0;
assign GPIO_2_OE_M2F[27:27]                           = GPIO_2_OE_M2F_net_1[27];
assign GPIO_2_OE_M2F_24_net_0[2]                      = GPIO_2_OE_M2F_24;
assign GPIO_2_OE_M2F[2:2]                             = GPIO_2_OE_M2F_24_net_0[2];
assign GPIO_2_OE_M2F_23_net_0[3]                      = GPIO_2_OE_M2F_23;
assign GPIO_2_OE_M2F[3:3]                             = GPIO_2_OE_M2F_23_net_0[3];
assign GPIO_2_OE_M2F_22_net_0[4]                      = GPIO_2_OE_M2F_22;
assign GPIO_2_OE_M2F[4:4]                             = GPIO_2_OE_M2F_22_net_0[4];
assign GPIO_2_OE_M2F_21_net_0[5]                      = GPIO_2_OE_M2F_21;
assign GPIO_2_OE_M2F[5:5]                             = GPIO_2_OE_M2F_21_net_0[5];
assign GPIO_2_OE_M2F_20_net_0[6]                      = GPIO_2_OE_M2F_20;
assign GPIO_2_OE_M2F[6:6]                             = GPIO_2_OE_M2F_20_net_0[6];
assign GPIO_2_OE_M2F_19_net_0[7]                      = GPIO_2_OE_M2F_19;
assign GPIO_2_OE_M2F[7:7]                             = GPIO_2_OE_M2F_19_net_0[7];
assign GPIO_2_OE_M2F_18_net_0[8]                      = GPIO_2_OE_M2F_18;
assign GPIO_2_OE_M2F[8:8]                             = GPIO_2_OE_M2F_18_net_0[8];
assign GPIO_2_OE_M2F_17_net_0[9]                      = GPIO_2_OE_M2F_17;
assign GPIO_2_OE_M2F[9:9]                             = GPIO_2_OE_M2F_17_net_0[9];
assign ADC_CSn_net_1                                  = ADC_CSn_net_0;
assign ADC_CSn                                        = ADC_CSn_net_1;
assign ADC_SCK_net_1                                  = ADC_SCK_net_0;
assign ADC_SCK                                        = ADC_SCK_net_1;
assign MMUART_2_TXD_net_1                             = MMUART_2_TXD_net_0;
assign MMUART_2_TXD                                   = MMUART_2_TXD_net_1;
assign MMUART_3_TXD_net_1                             = MMUART_3_TXD_net_0;
assign MMUART_3_TXD                                   = MMUART_3_TXD_net_1;
assign MMUART_4_TXD_net_1                             = MMUART_4_TXD_net_0;
assign MMUART_4_TXD                                   = MMUART_4_TXD_net_1;
assign PHY_MDC_net_1                                  = PHY_MDC_net_0;
assign PHY_MDC                                        = PHY_MDC_net_1;
assign M2_W_DISABLE1_net_1                            = M2_W_DISABLE1_net_0;
assign M2_W_DISABLE1                                  = M2_W_DISABLE1_net_1;
assign M2_W_DISABLE2_net_1                            = M2_W_DISABLE2_net_0;
assign M2_W_DISABLE2                                  = M2_W_DISABLE2_net_1;
assign MAC_1_MDO_OE_M2F_net_1                         = MAC_1_MDO_OE_M2F_net_0;
assign MAC_1_MDO_OE_M2F                               = MAC_1_MDO_OE_M2F_net_1;
assign MAC_1_MDC_M2F_net_1                            = MAC_1_MDC_M2F_net_0;
assign MAC_1_MDC_M2F                                  = MAC_1_MDC_M2F_net_1;
assign MAC_1_MDO_M2F_net_1                            = MAC_1_MDO_M2F_net_0;
assign MAC_1_MDO_M2F                                  = MAC_1_MDO_M2F_net_1;
assign EMMC_CLK_net_1                                 = EMMC_CLK_net_0;
assign EMMC_CLK                                       = EMMC_CLK_net_1;
assign EMMC_RSTN_net_1                                = EMMC_RSTN_net_0;
assign EMMC_RSTN                                      = EMMC_RSTN_net_1;
assign VIO_ENABLE_net_1                               = VIO_ENABLE_net_0;
assign VIO_ENABLE                                     = VIO_ENABLE_net_1;
assign FIC_2_AXI4_TARGET_AWREADY_net_0                = FIC_2_AXI4_TARGET_AWREADY;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWREADY         = FIC_2_AXI4_TARGET_AWREADY_net_0;
assign FIC_2_AXI4_TARGET_WREADY_net_0                 = FIC_2_AXI4_TARGET_WREADY;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WREADY          = FIC_2_AXI4_TARGET_WREADY_net_0;
assign FIC_2_AXI4_TARGET_BID_net_0                    = FIC_2_AXI4_TARGET_BID;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BID[3:0]        = FIC_2_AXI4_TARGET_BID_net_0;
assign FIC_2_AXI4_TARGET_BRESP_net_0                  = FIC_2_AXI4_TARGET_BRESP;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BRESP[1:0]      = FIC_2_AXI4_TARGET_BRESP_net_0;
assign FIC_2_AXI4_TARGET_BVALID_net_0                 = FIC_2_AXI4_TARGET_BVALID;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BVALID          = FIC_2_AXI4_TARGET_BVALID_net_0;
assign FIC_2_AXI4_TARGET_ARREADY_net_0                = FIC_2_AXI4_TARGET_ARREADY;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARREADY         = FIC_2_AXI4_TARGET_ARREADY_net_0;
assign FIC_2_AXI4_TARGET_RID_net_0                    = FIC_2_AXI4_TARGET_RID;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RID[3:0]        = FIC_2_AXI4_TARGET_RID_net_0;
assign FIC_2_AXI4_TARGET_RDATA_net_0                  = FIC_2_AXI4_TARGET_RDATA;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RDATA[63:0]     = FIC_2_AXI4_TARGET_RDATA_net_0;
assign FIC_2_AXI4_TARGET_RRESP_net_0                  = FIC_2_AXI4_TARGET_RRESP;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RRESP[1:0]      = FIC_2_AXI4_TARGET_RRESP_net_0;
assign FIC_2_AXI4_TARGET_RLAST_net_0                  = FIC_2_AXI4_TARGET_RLAST;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RLAST           = FIC_2_AXI4_TARGET_RLAST_net_0;
assign FIC_2_AXI4_TARGET_RVALID_net_0                 = FIC_2_AXI4_TARGET_RVALID;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RVALID          = FIC_2_AXI4_TARGET_RVALID_net_0;
assign FIC_1_AXI4_TARGET_AWREADY_net_0                = FIC_1_AXI4_TARGET_AWREADY;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWREADY         = FIC_1_AXI4_TARGET_AWREADY_net_0;
assign FIC_1_AXI4_TARGET_WREADY_net_0                 = FIC_1_AXI4_TARGET_WREADY;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WREADY          = FIC_1_AXI4_TARGET_WREADY_net_0;
assign FIC_1_AXI4_TARGET_BID_net_0                    = FIC_1_AXI4_TARGET_BID;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BID[3:0]        = FIC_1_AXI4_TARGET_BID_net_0;
assign FIC_1_AXI4_TARGET_BRESP_net_0                  = FIC_1_AXI4_TARGET_BRESP;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BRESP[1:0]      = FIC_1_AXI4_TARGET_BRESP_net_0;
assign FIC_1_AXI4_TARGET_BVALID_net_0                 = FIC_1_AXI4_TARGET_BVALID;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BVALID          = FIC_1_AXI4_TARGET_BVALID_net_0;
assign FIC_1_AXI4_TARGET_ARREADY_net_0                = FIC_1_AXI4_TARGET_ARREADY;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARREADY         = FIC_1_AXI4_TARGET_ARREADY_net_0;
assign FIC_1_AXI4_TARGET_RID_net_0                    = FIC_1_AXI4_TARGET_RID;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RID[3:0]        = FIC_1_AXI4_TARGET_RID_net_0;
assign FIC_1_AXI4_TARGET_RDATA_net_0                  = FIC_1_AXI4_TARGET_RDATA;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RDATA[63:0]     = FIC_1_AXI4_TARGET_RDATA_net_0;
assign FIC_1_AXI4_TARGET_RRESP_net_0                  = FIC_1_AXI4_TARGET_RRESP;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RRESP[1:0]      = FIC_1_AXI4_TARGET_RRESP_net_0;
assign FIC_1_AXI4_TARGET_RLAST_net_0                  = FIC_1_AXI4_TARGET_RLAST;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RLAST           = FIC_1_AXI4_TARGET_RLAST_net_0;
assign FIC_1_AXI4_TARGET_RVALID_net_0                 = FIC_1_AXI4_TARGET_RVALID;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RVALID          = FIC_1_AXI4_TARGET_RVALID_net_0;
assign FIC_0_AXI4_TARGET_AWREADY_net_0                = FIC_0_AXI4_TARGET_AWREADY;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWREADY         = FIC_0_AXI4_TARGET_AWREADY_net_0;
assign FIC_0_AXI4_TARGET_WREADY_net_0                 = FIC_0_AXI4_TARGET_WREADY;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WREADY          = FIC_0_AXI4_TARGET_WREADY_net_0;
assign FIC_0_AXI4_TARGET_BID_net_0                    = FIC_0_AXI4_TARGET_BID;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BID[3:0]        = FIC_0_AXI4_TARGET_BID_net_0;
assign FIC_0_AXI4_TARGET_BRESP_net_0                  = FIC_0_AXI4_TARGET_BRESP;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BRESP[1:0]      = FIC_0_AXI4_TARGET_BRESP_net_0;
assign FIC_0_AXI4_TARGET_BVALID_net_0                 = FIC_0_AXI4_TARGET_BVALID;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BVALID          = FIC_0_AXI4_TARGET_BVALID_net_0;
assign FIC_0_AXI4_TARGET_ARREADY_net_0                = FIC_0_AXI4_TARGET_ARREADY;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARREADY         = FIC_0_AXI4_TARGET_ARREADY_net_0;
assign FIC_0_AXI4_TARGET_RID_net_0                    = FIC_0_AXI4_TARGET_RID;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RID[3:0]        = FIC_0_AXI4_TARGET_RID_net_0;
assign FIC_0_AXI4_TARGET_RDATA_net_0                  = FIC_0_AXI4_TARGET_RDATA;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RDATA[63:0]     = FIC_0_AXI4_TARGET_RDATA_net_0;
assign FIC_0_AXI4_TARGET_RRESP_net_0                  = FIC_0_AXI4_TARGET_RRESP;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RRESP[1:0]      = FIC_0_AXI4_TARGET_RRESP_net_0;
assign FIC_0_AXI4_TARGET_RLAST_net_0                  = FIC_0_AXI4_TARGET_RLAST;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RLAST           = FIC_0_AXI4_TARGET_RLAST_net_0;
assign FIC_0_AXI4_TARGET_RVALID_net_0                 = FIC_0_AXI4_TARGET_RVALID;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RVALID          = FIC_0_AXI4_TARGET_RVALID_net_0;
assign CAPE_APB_MTARGET_PADDR_net_0                   = CAPE_APB_MTARGET_PADDR;
assign CAPE_APB_MTARGET_PADDRS[31:0]                  = CAPE_APB_MTARGET_PADDR_net_0;
assign CAPE_APB_MTARGET_PSELx_net_0                   = CAPE_APB_MTARGET_PSELx;
assign CAPE_APB_MTARGET_PSELS1                        = CAPE_APB_MTARGET_PSELx_net_0;
assign CAPE_APB_MTARGET_PENABLE_net_0                 = CAPE_APB_MTARGET_PENABLE;
assign CAPE_APB_MTARGET_PENABLES                      = CAPE_APB_MTARGET_PENABLE_net_0;
assign CAPE_APB_MTARGET_PWRITE_net_0                  = CAPE_APB_MTARGET_PWRITE;
assign CAPE_APB_MTARGET_PWRITES                       = CAPE_APB_MTARGET_PWRITE_net_0;
assign CAPE_APB_MTARGET_PWDATA_net_0                  = CAPE_APB_MTARGET_PWDATA;
assign CAPE_APB_MTARGET_PWDATAS[31:0]                 = CAPE_APB_MTARGET_PWDATA_net_0;
assign CSI_APB_MTARGET_PSELx_net_0                    = CSI_APB_MTARGET_PSELx;
assign CSI_APB_MTARGET_PSELS2                         = CSI_APB_MTARGET_PSELx_net_0;
assign HSI_APB_MTARGET_PSELx_net_0                    = HSI_APB_MTARGET_PSELx;
assign HSI_APB_MTARGET_PSELS4                         = HSI_APB_MTARGET_PSELx_net_0;
assign M2_APB_MTARGET_PSELx_net_0                     = M2_APB_MTARGET_PSELx;
assign M2_APB_MTARGET_PSELS16                         = M2_APB_MTARGET_PSELx_net_0;
assign MSS_RESET_N_M2F_net_1                          = MSS_RESET_N_M2F_net_0;
assign MSS_RESET_N_M2F                                = MSS_RESET_N_M2F_net_1;
assign FIC_3_APB_M_PSTRB_net_1                        = FIC_3_APB_M_PSTRB_net_0;
assign FIC_3_APB_M_PSTRB[3:0]                         = FIC_3_APB_M_PSTRB_net_1;
assign FIC_0_AXI4_INITIATOR_AWID_net_0                = FIC_0_AXI4_INITIATOR_AWID;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWID[7:0]    = FIC_0_AXI4_INITIATOR_AWID_net_0;
assign FIC_0_AXI4_INITIATOR_AWADDR_net_0              = FIC_0_AXI4_INITIATOR_AWADDR;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWADDR[37:0] = FIC_0_AXI4_INITIATOR_AWADDR_net_0;
assign FIC_0_AXI4_INITIATOR_AWLEN_net_0               = FIC_0_AXI4_INITIATOR_AWLEN;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWLEN[7:0]   = FIC_0_AXI4_INITIATOR_AWLEN_net_0;
assign FIC_0_AXI4_INITIATOR_AWSIZE_net_0              = FIC_0_AXI4_INITIATOR_AWSIZE;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWSIZE[2:0]  = FIC_0_AXI4_INITIATOR_AWSIZE_net_0;
assign FIC_0_AXI4_INITIATOR_AWBURST_net_0             = FIC_0_AXI4_INITIATOR_AWBURST;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWBURST[1:0] = FIC_0_AXI4_INITIATOR_AWBURST_net_0;
assign FIC_0_AXI4_INITIATOR_AWLOCK_net_0              = FIC_0_AXI4_INITIATOR_AWLOCK;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWLOCK       = FIC_0_AXI4_INITIATOR_AWLOCK_net_0;
assign FIC_0_AXI4_INITIATOR_AWQOS_net_0               = FIC_0_AXI4_INITIATOR_AWQOS;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWQOS[3:0]   = FIC_0_AXI4_INITIATOR_AWQOS_net_0;
assign FIC_0_AXI4_INITIATOR_AWCACHE_net_0             = FIC_0_AXI4_INITIATOR_AWCACHE;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWCACHE[3:0] = FIC_0_AXI4_INITIATOR_AWCACHE_net_0;
assign FIC_0_AXI4_INITIATOR_AWPROT_net_0              = FIC_0_AXI4_INITIATOR_AWPROT;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWPROT[2:0]  = FIC_0_AXI4_INITIATOR_AWPROT_net_0;
assign FIC_0_AXI4_INITIATOR_AWVALID_net_0             = FIC_0_AXI4_INITIATOR_AWVALID;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWVALID      = FIC_0_AXI4_INITIATOR_AWVALID_net_0;
assign FIC_0_AXI4_INITIATOR_WDATA_net_0               = FIC_0_AXI4_INITIATOR_WDATA;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WDATA[63:0]  = FIC_0_AXI4_INITIATOR_WDATA_net_0;
assign FIC_0_AXI4_INITIATOR_WSTRB_net_0               = FIC_0_AXI4_INITIATOR_WSTRB;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WSTRB[7:0]   = FIC_0_AXI4_INITIATOR_WSTRB_net_0;
assign FIC_0_AXI4_INITIATOR_WLAST_net_0               = FIC_0_AXI4_INITIATOR_WLAST;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WLAST        = FIC_0_AXI4_INITIATOR_WLAST_net_0;
assign FIC_0_AXI4_INITIATOR_WVALID_net_0              = FIC_0_AXI4_INITIATOR_WVALID;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WVALID       = FIC_0_AXI4_INITIATOR_WVALID_net_0;
assign FIC_0_AXI4_INITIATOR_BREADY_net_0              = FIC_0_AXI4_INITIATOR_BREADY;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BREADY       = FIC_0_AXI4_INITIATOR_BREADY_net_0;
assign FIC_0_AXI4_INITIATOR_ARID_net_0                = FIC_0_AXI4_INITIATOR_ARID;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARID[7:0]    = FIC_0_AXI4_INITIATOR_ARID_net_0;
assign FIC_0_AXI4_INITIATOR_ARADDR_net_0              = FIC_0_AXI4_INITIATOR_ARADDR;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARADDR[37:0] = FIC_0_AXI4_INITIATOR_ARADDR_net_0;
assign FIC_0_AXI4_INITIATOR_ARLEN_net_0               = FIC_0_AXI4_INITIATOR_ARLEN;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARLEN[7:0]   = FIC_0_AXI4_INITIATOR_ARLEN_net_0;
assign FIC_0_AXI4_INITIATOR_ARSIZE_net_0              = FIC_0_AXI4_INITIATOR_ARSIZE;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARSIZE[2:0]  = FIC_0_AXI4_INITIATOR_ARSIZE_net_0;
assign FIC_0_AXI4_INITIATOR_ARBURST_net_0             = FIC_0_AXI4_INITIATOR_ARBURST;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARBURST[1:0] = FIC_0_AXI4_INITIATOR_ARBURST_net_0;
assign FIC_0_AXI4_INITIATOR_ARLOCK_net_0              = FIC_0_AXI4_INITIATOR_ARLOCK;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARLOCK       = FIC_0_AXI4_INITIATOR_ARLOCK_net_0;
assign FIC_0_AXI4_INITIATOR_ARQOS_net_0               = FIC_0_AXI4_INITIATOR_ARQOS;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARQOS[3:0]   = FIC_0_AXI4_INITIATOR_ARQOS_net_0;
assign FIC_0_AXI4_INITIATOR_ARCACHE_net_0             = FIC_0_AXI4_INITIATOR_ARCACHE;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARCACHE[3:0] = FIC_0_AXI4_INITIATOR_ARCACHE_net_0;
assign FIC_0_AXI4_INITIATOR_ARPROT_net_0              = FIC_0_AXI4_INITIATOR_ARPROT;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARPROT[2:0]  = FIC_0_AXI4_INITIATOR_ARPROT_net_0;
assign FIC_0_AXI4_INITIATOR_ARVALID_net_0             = FIC_0_AXI4_INITIATOR_ARVALID;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARVALID      = FIC_0_AXI4_INITIATOR_ARVALID_net_0;
assign FIC_0_AXI4_INITIATOR_RREADY_net_0              = FIC_0_AXI4_INITIATOR_RREADY;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RREADY       = FIC_0_AXI4_INITIATOR_RREADY_net_0;
assign FIC_1_AXI4_INITIATOR_AWID_net_0                = FIC_1_AXI4_INITIATOR_AWID;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWID[7:0]    = FIC_1_AXI4_INITIATOR_AWID_net_0;
assign FIC_1_AXI4_INITIATOR_AWADDR_net_0              = FIC_1_AXI4_INITIATOR_AWADDR;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWADDR[37:0] = FIC_1_AXI4_INITIATOR_AWADDR_net_0;
assign FIC_1_AXI4_INITIATOR_AWLEN_net_0               = FIC_1_AXI4_INITIATOR_AWLEN;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWLEN[7:0]   = FIC_1_AXI4_INITIATOR_AWLEN_net_0;
assign FIC_1_AXI4_INITIATOR_AWSIZE_net_0              = FIC_1_AXI4_INITIATOR_AWSIZE;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWSIZE[2:0]  = FIC_1_AXI4_INITIATOR_AWSIZE_net_0;
assign FIC_1_AXI4_INITIATOR_AWBURST_net_0             = FIC_1_AXI4_INITIATOR_AWBURST;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWBURST[1:0] = FIC_1_AXI4_INITIATOR_AWBURST_net_0;
assign FIC_1_AXI4_INITIATOR_AWLOCK_net_0              = FIC_1_AXI4_INITIATOR_AWLOCK;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWLOCK       = FIC_1_AXI4_INITIATOR_AWLOCK_net_0;
assign FIC_1_AXI4_INITIATOR_AWQOS_net_0               = FIC_1_AXI4_INITIATOR_AWQOS;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWQOS[3:0]   = FIC_1_AXI4_INITIATOR_AWQOS_net_0;
assign FIC_1_AXI4_INITIATOR_AWCACHE_net_0             = FIC_1_AXI4_INITIATOR_AWCACHE;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWCACHE[3:0] = FIC_1_AXI4_INITIATOR_AWCACHE_net_0;
assign FIC_1_AXI4_INITIATOR_AWPROT_net_0              = FIC_1_AXI4_INITIATOR_AWPROT;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWPROT[2:0]  = FIC_1_AXI4_INITIATOR_AWPROT_net_0;
assign FIC_1_AXI4_INITIATOR_AWVALID_net_0             = FIC_1_AXI4_INITIATOR_AWVALID;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWVALID      = FIC_1_AXI4_INITIATOR_AWVALID_net_0;
assign FIC_1_AXI4_INITIATOR_WDATA_net_0               = FIC_1_AXI4_INITIATOR_WDATA;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WDATA[63:0]  = FIC_1_AXI4_INITIATOR_WDATA_net_0;
assign FIC_1_AXI4_INITIATOR_WSTRB_net_0               = FIC_1_AXI4_INITIATOR_WSTRB;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WSTRB[7:0]   = FIC_1_AXI4_INITIATOR_WSTRB_net_0;
assign FIC_1_AXI4_INITIATOR_WLAST_net_0               = FIC_1_AXI4_INITIATOR_WLAST;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WLAST        = FIC_1_AXI4_INITIATOR_WLAST_net_0;
assign FIC_1_AXI4_INITIATOR_WVALID_net_0              = FIC_1_AXI4_INITIATOR_WVALID;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WVALID       = FIC_1_AXI4_INITIATOR_WVALID_net_0;
assign FIC_1_AXI4_INITIATOR_BREADY_net_0              = FIC_1_AXI4_INITIATOR_BREADY;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BREADY       = FIC_1_AXI4_INITIATOR_BREADY_net_0;
assign FIC_1_AXI4_INITIATOR_ARID_net_0                = FIC_1_AXI4_INITIATOR_ARID;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARID[7:0]    = FIC_1_AXI4_INITIATOR_ARID_net_0;
assign FIC_1_AXI4_INITIATOR_ARADDR_net_0              = FIC_1_AXI4_INITIATOR_ARADDR;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARADDR[37:0] = FIC_1_AXI4_INITIATOR_ARADDR_net_0;
assign FIC_1_AXI4_INITIATOR_ARLEN_net_0               = FIC_1_AXI4_INITIATOR_ARLEN;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARLEN[7:0]   = FIC_1_AXI4_INITIATOR_ARLEN_net_0;
assign FIC_1_AXI4_INITIATOR_ARSIZE_net_0              = FIC_1_AXI4_INITIATOR_ARSIZE;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARSIZE[2:0]  = FIC_1_AXI4_INITIATOR_ARSIZE_net_0;
assign FIC_1_AXI4_INITIATOR_ARBURST_net_0             = FIC_1_AXI4_INITIATOR_ARBURST;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARBURST[1:0] = FIC_1_AXI4_INITIATOR_ARBURST_net_0;
assign FIC_1_AXI4_INITIATOR_ARLOCK_net_0              = FIC_1_AXI4_INITIATOR_ARLOCK;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARLOCK       = FIC_1_AXI4_INITIATOR_ARLOCK_net_0;
assign FIC_1_AXI4_INITIATOR_ARQOS_net_0               = FIC_1_AXI4_INITIATOR_ARQOS;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARQOS[3:0]   = FIC_1_AXI4_INITIATOR_ARQOS_net_0;
assign FIC_1_AXI4_INITIATOR_ARCACHE_net_0             = FIC_1_AXI4_INITIATOR_ARCACHE;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARCACHE[3:0] = FIC_1_AXI4_INITIATOR_ARCACHE_net_0;
assign FIC_1_AXI4_INITIATOR_ARPROT_net_0              = FIC_1_AXI4_INITIATOR_ARPROT;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARPROT[2:0]  = FIC_1_AXI4_INITIATOR_ARPROT_net_0;
assign FIC_1_AXI4_INITIATOR_ARVALID_net_0             = FIC_1_AXI4_INITIATOR_ARVALID;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARVALID      = FIC_1_AXI4_INITIATOR_ARVALID_net_0;
assign FIC_1_AXI4_INITIATOR_RREADY_net_0              = FIC_1_AXI4_INITIATOR_RREADY;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RREADY       = FIC_1_AXI4_INITIATOR_RREADY_net_0;
assign SPI_0_CLK_net_1                                = SPI_0_CLK_net_0;
assign SPI_0_CLK                                      = SPI_0_CLK_net_1;
assign SPI_0_DO_net_1                                 = SPI_0_DO_net_0;
assign SPI_0_DO                                       = SPI_0_DO_net_1;
assign SPI_0_SS1_net_1                                = SPI_0_SS1_net_0;
assign SPI_0_SS1                                      = SPI_0_SS1_net_1;
assign SPI_1_SS1_net_1                                = SPI_1_SS1_net_0;
assign SPI_1_SS1                                      = SPI_1_SS1_net_1;
assign SPI_1_CLK_net_1                                = SPI_1_CLK_net_0;
assign SPI_1_CLK                                      = SPI_1_CLK_net_1;
assign SPI_1_DO_net_1                                 = SPI_1_DO_net_0;
assign SPI_1_DO                                       = SPI_1_DO_net_1;
//--------------------------------------------------------------------
// Slices assignments
//--------------------------------------------------------------------
assign GPIO_2_F2M_slice_0[27]  = GPIO_2_F2M[27:27];
assign GPIO_2_F2M_slice_1[26]  = GPIO_2_F2M[26:26];
assign GPIO_2_F2M_slice_2[25]  = GPIO_2_F2M[25:25];
assign GPIO_2_F2M_slice_3[24]  = GPIO_2_F2M[24:24];
assign GPIO_2_F2M_slice_4[23]  = GPIO_2_F2M[23:23];
assign GPIO_2_F2M_slice_5[22]  = GPIO_2_F2M[22:22];
assign GPIO_2_F2M_slice_6[21]  = GPIO_2_F2M[21:21];
assign GPIO_2_F2M_slice_7[20]  = GPIO_2_F2M[20:20];
assign GPIO_2_F2M_slice_8[19]  = GPIO_2_F2M[19:19];
assign GPIO_2_F2M_slice_9[18]  = GPIO_2_F2M[18:18];
assign GPIO_2_F2M_slice_10[17] = GPIO_2_F2M[17:17];
assign GPIO_2_F2M_slice_11[16] = GPIO_2_F2M[16:16];
assign GPIO_2_F2M_slice_12[15] = GPIO_2_F2M[15:15];
assign GPIO_2_F2M_slice_13[14] = GPIO_2_F2M[14:14];
assign GPIO_2_F2M_slice_14[13] = GPIO_2_F2M[13:13];
assign GPIO_2_F2M_slice_15[12] = GPIO_2_F2M[12:12];
assign GPIO_2_F2M_slice_16[11] = GPIO_2_F2M[11:11];
assign GPIO_2_F2M_slice_17[10] = GPIO_2_F2M[10:10];
assign GPIO_2_F2M_slice_18[9]  = GPIO_2_F2M[9:9];
assign GPIO_2_F2M_slice_19[8]  = GPIO_2_F2M[8:8];
assign GPIO_2_F2M_slice_20[7]  = GPIO_2_F2M[7:7];
assign GPIO_2_F2M_slice_21[6]  = GPIO_2_F2M[6:6];
assign GPIO_2_F2M_slice_22[5]  = GPIO_2_F2M[5:5];
assign GPIO_2_F2M_slice_23[4]  = GPIO_2_F2M[4:4];
assign GPIO_2_F2M_slice_24[3]  = GPIO_2_F2M[3:3];
assign GPIO_2_F2M_slice_25[2]  = GPIO_2_F2M[2:2];
assign GPIO_2_F2M_slice_26[1]  = GPIO_2_F2M[1:1];
assign GPIO_2_F2M_slice_27[0]  = GPIO_2_F2M[0:0];
//--------------------------------------------------------------------
// Concatenation assignments
//--------------------------------------------------------------------
assign MSS_INT_F2M_net_0 = { IHC_SUBSYSTEM_0_E51_IRQ , IHC_SUBSYSTEM_0_U54_1_IRQ , IHC_SUBSYSTEM_0_U54_2_IRQ , IHC_SUBSYSTEM_0_U54_3_IRQ , IHC_SUBSYSTEM_0_U54_4_IRQ , MSS_INT_F2M , PHY_INTn , PCIE_INT , 1'b0 };
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------AND4
AND4 AND_DLL_LOCKS(
        // Inputs
        .A ( PF_SOC_MSS_FIC_0_DLL_LOCK_M2F ),
        .B ( PF_SOC_MSS_FIC_1_DLL_LOCK_M2F ),
        .C ( PF_SOC_MSS_FIC_2_DLL_LOCK_M2F ),
        .D ( PF_SOC_MSS_FIC_3_DLL_LOCK_M2F ),
        // Outputs
        .Y ( MSS_DLL_LOCKS_net_0 ) 
        );

//--------APB_ARBITER
APB_ARBITER #( 
        .select_bit ( 28 ) )
APB_ARBITER_0(
        // Inputs
        .in_penable       ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PENABLE ),
        .in_psel          ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PSELx ),
        .in_paddr         ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PADDR ),
        .in_pwrite        ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PWRITE ),
        .in_pwdata        ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PWDATA ),
        .out_low_prdata   ( APB_ARBITER_0_APB_MASTER_low_PRDATA ),
        .out_low_pready   ( APB_ARBITER_0_APB_MASTER_low_PREADY ),
        .out_low_pslverr  ( APB_ARBITER_0_APB_MASTER_low_PSLVERR ),
        .out_high_prdata  ( APB_ARBITER_0_APB_MASTER_high_PRDATA ),
        .out_high_pready  ( APB_ARBITER_0_APB_MASTER_high_PREADY ),
        .out_high_pslverr ( APB_ARBITER_0_APB_MASTER_high_PSLVERR ),
        // Outputs
        .in_prdata        ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PRDATA ),
        .in_pready        ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PREADY ),
        .in_pslverr       ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PSLVERR ),
        .out_low_penable  ( APB_ARBITER_0_APB_MASTER_low_PENABLE ),
        .out_low_psel     ( APB_ARBITER_0_APB_MASTER_low_PSELx ),
        .out_low_paddr    ( APB_ARBITER_0_APB_MASTER_low_PADDR ),
        .out_low_pwrite   ( APB_ARBITER_0_APB_MASTER_low_PWRITE ),
        .out_low_pwdata   ( APB_ARBITER_0_APB_MASTER_low_PWDATA ),
        .out_high_penable ( APB_ARBITER_0_APB_MASTER_high_PENABLE ),
        .out_high_psel    ( APB_ARBITER_0_APB_MASTER_high_PSELx ),
        .out_high_paddr   ( APB_ARBITER_0_APB_MASTER_high_PADDR ),
        .out_high_pwrite  ( APB_ARBITER_0_APB_MASTER_high_PWRITE ),
        .out_high_pwdata  ( APB_ARBITER_0_APB_MASTER_high_PWDATA ) 
        );

//--------FIC3_INITIATOR
FIC3_INITIATOR FIC3_INITIATOR_inst_0(
        // Inputs
        .PADDR      ( APB_ARBITER_0_APB_MASTER_low_PADDR ),
        .PSEL       ( APB_ARBITER_0_APB_MASTER_low_PSELx ),
        .PENABLE    ( APB_ARBITER_0_APB_MASTER_low_PENABLE ),
        .PWRITE     ( APB_ARBITER_0_APB_MASTER_low_PWRITE ),
        .PWDATA     ( APB_ARBITER_0_APB_MASTER_low_PWDATA ),
        .PRDATAS1   ( CAPE_APB_MTARGET_PRDATAS1 ),
        .PREADYS1   ( CAPE_APB_MTARGET_PREADYS1 ),
        .PSLVERRS1  ( CAPE_APB_MTARGET_PSLVERRS1 ),
        .PRDATAS2   ( CSI_APB_MTARGET_PRDATAS2 ),
        .PREADYS2   ( CSI_APB_MTARGET_PREADYS2 ),
        .PSLVERRS2  ( CSI_APB_MTARGET_PSLVERRS2 ),
        .PRDATAS4   ( HSI_APB_MTARGET_PRDATAS4 ),
        .PREADYS4   ( HSI_APB_MTARGET_PREADYS4 ),
        .PSLVERRS4  ( HSI_APB_MTARGET_PSLVERRS4 ),
        .PRDATAS16  ( M2_APB_MTARGET_PRDATAS16 ),
        .PREADYS16  ( M2_APB_MTARGET_PREADYS16 ),
        .PSLVERRS16 ( M2_APB_MTARGET_PSLVERRS16 ),
        // Outputs
        .PRDATA     ( APB_ARBITER_0_APB_MASTER_low_PRDATA ),
        .PREADY     ( APB_ARBITER_0_APB_MASTER_low_PREADY ),
        .PSLVERR    ( APB_ARBITER_0_APB_MASTER_low_PSLVERR ),
        .PADDRS     ( CAPE_APB_MTARGET_PADDR ),
        .PSELS1     ( CAPE_APB_MTARGET_PSELx ),
        .PENABLES   ( CAPE_APB_MTARGET_PENABLE ),
        .PWRITES    ( CAPE_APB_MTARGET_PWRITE ),
        .PWDATAS    ( CAPE_APB_MTARGET_PWDATA ),
        .PSELS2     ( CSI_APB_MTARGET_PSELx ),
        .PSELS4     ( HSI_APB_MTARGET_PSELx ),
        .PSELS16    ( M2_APB_MTARGET_PSELx ) 
        );

//--------BIBUF
BIBUF I2C0_SCL_BIBUF(
        // Inputs
        .D   ( GND_net ),
        .E   ( PF_SOC_MSS_I2C_0_SCL_OE_M2F ),
        // Outputs
        .Y   ( I2C0_SCL_BIBUF_Y ),
        // Inouts
        .PAD ( I2C0_SCL ) 
        );

//--------BIBUF
BIBUF I2C0_SDA_BIBUF(
        // Inputs
        .D   ( GND_net ),
        .E   ( PF_SOC_MSS_I2C_0_SDA_OE_M2F ),
        // Outputs
        .Y   ( I2C0_SDA_BIBUF_Y ),
        // Inouts
        .PAD ( I2C0_SDA ) 
        );

//--------IHC_SUBSYSTEM
IHC_SUBSYSTEM IHC_SUBSYSTEM_0(
        // Inputs
        .presetn   ( PRESETN ),
        .pclk      ( FIC_3_PCLK ),
        .PSEL      ( APB_ARBITER_0_APB_MASTER_high_PSELx ),
        .PENABLE   ( APB_ARBITER_0_APB_MASTER_high_PENABLE ),
        .PWRITE    ( APB_ARBITER_0_APB_MASTER_high_PWRITE ),
        .PADDR     ( APB_ARBITER_0_APB_MASTER_high_PADDR ),
        .PWDATA    ( APB_ARBITER_0_APB_MASTER_high_PWDATA ),
        // Outputs
        .E51_IRQ   ( IHC_SUBSYSTEM_0_E51_IRQ ),
        .PREADY    ( APB_ARBITER_0_APB_MASTER_high_PREADY ),
        .PSLVERR   ( APB_ARBITER_0_APB_MASTER_high_PSLVERR ),
        .U54_1_IRQ ( IHC_SUBSYSTEM_0_U54_1_IRQ ),
        .U54_2_IRQ ( IHC_SUBSYSTEM_0_U54_2_IRQ ),
        .U54_3_IRQ ( IHC_SUBSYSTEM_0_U54_3_IRQ ),
        .U54_4_IRQ ( IHC_SUBSYSTEM_0_U54_4_IRQ ),
        .PRDATA    ( APB_ARBITER_0_APB_MASTER_high_PRDATA ) 
        );

//--------PF_SOC_MSS
PF_SOC_MSS PF_SOC_MSS_inst_0(
        // Inputs
        .FIC_0_ACLK           ( FIC_0_ACLK ),
        .FIC_0_AXI4_M_AWREADY ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWREADY ),
        .FIC_0_AXI4_M_WREADY  ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WREADY ),
        .FIC_0_AXI4_M_BID     ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BID ),
        .FIC_0_AXI4_M_BRESP   ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BRESP ),
        .FIC_0_AXI4_M_BVALID  ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BVALID ),
        .FIC_0_AXI4_M_ARREADY ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARREADY ),
        .FIC_0_AXI4_M_RID     ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RID ),
        .FIC_0_AXI4_M_RDATA   ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RDATA ),
        .FIC_0_AXI4_M_RRESP   ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RRESP ),
        .FIC_0_AXI4_M_RLAST   ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RLAST ),
        .FIC_0_AXI4_M_RVALID  ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RVALID ),
        .FIC_0_AXI4_S_AWID    ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWID ),
        .FIC_0_AXI4_S_AWADDR  ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWADDR ),
        .FIC_0_AXI4_S_AWLEN   ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLEN ),
        .FIC_0_AXI4_S_AWSIZE  ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWSIZE ),
        .FIC_0_AXI4_S_AWBURST ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWBURST ),
        .FIC_0_AXI4_S_AWQOS   ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWQOS ),
        .FIC_0_AXI4_S_AWLOCK  ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLOCK ),
        .FIC_0_AXI4_S_AWCACHE ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWCACHE ),
        .FIC_0_AXI4_S_AWPROT  ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWPROT ),
        .FIC_0_AXI4_S_AWVALID ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWVALID ),
        .FIC_0_AXI4_S_WDATA   ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WDATA ),
        .FIC_0_AXI4_S_WSTRB   ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WSTRB ),
        .FIC_0_AXI4_S_WLAST   ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WLAST ),
        .FIC_0_AXI4_S_WVALID  ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WVALID ),
        .FIC_0_AXI4_S_BREADY  ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BREADY ),
        .FIC_0_AXI4_S_ARID    ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARID ),
        .FIC_0_AXI4_S_ARADDR  ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARADDR ),
        .FIC_0_AXI4_S_ARLEN   ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLEN ),
        .FIC_0_AXI4_S_ARSIZE  ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARSIZE ),
        .FIC_0_AXI4_S_ARBURST ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARBURST ),
        .FIC_0_AXI4_S_ARQOS   ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARQOS ),
        .FIC_0_AXI4_S_ARLOCK  ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLOCK ),
        .FIC_0_AXI4_S_ARCACHE ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARCACHE ),
        .FIC_0_AXI4_S_ARPROT  ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARPROT ),
        .FIC_0_AXI4_S_ARVALID ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARVALID ),
        .FIC_0_AXI4_S_RREADY  ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RREADY ),
        .FIC_1_ACLK           ( FIC_1_ACLK ),
        .FIC_1_AXI4_M_AWREADY ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWREADY ),
        .FIC_1_AXI4_M_WREADY  ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WREADY ),
        .FIC_1_AXI4_M_BID     ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BID ),
        .FIC_1_AXI4_M_BRESP   ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BRESP ),
        .FIC_1_AXI4_M_BVALID  ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BVALID ),
        .FIC_1_AXI4_M_ARREADY ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARREADY ),
        .FIC_1_AXI4_M_RID     ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RID ),
        .FIC_1_AXI4_M_RDATA   ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RDATA ),
        .FIC_1_AXI4_M_RRESP   ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RRESP ),
        .FIC_1_AXI4_M_RLAST   ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RLAST ),
        .FIC_1_AXI4_M_RVALID  ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RVALID ),
        .FIC_1_AXI4_S_AWID    ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWID ),
        .FIC_1_AXI4_S_AWADDR  ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWADDR ),
        .FIC_1_AXI4_S_AWLEN   ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLEN ),
        .FIC_1_AXI4_S_AWSIZE  ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWSIZE ),
        .FIC_1_AXI4_S_AWBURST ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWBURST ),
        .FIC_1_AXI4_S_AWLOCK  ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLOCK ),
        .FIC_1_AXI4_S_AWCACHE ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWCACHE ),
        .FIC_1_AXI4_S_AWQOS   ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWQOS ),
        .FIC_1_AXI4_S_AWPROT  ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWPROT ),
        .FIC_1_AXI4_S_AWVALID ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWVALID ),
        .FIC_1_AXI4_S_WDATA   ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WDATA ),
        .FIC_1_AXI4_S_WSTRB   ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WSTRB ),
        .FIC_1_AXI4_S_WLAST   ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WLAST ),
        .FIC_1_AXI4_S_WVALID  ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WVALID ),
        .FIC_1_AXI4_S_BREADY  ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BREADY ),
        .FIC_1_AXI4_S_ARID    ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARID ),
        .FIC_1_AXI4_S_ARADDR  ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARADDR ),
        .FIC_1_AXI4_S_ARLEN   ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLEN ),
        .FIC_1_AXI4_S_ARSIZE  ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARSIZE ),
        .FIC_1_AXI4_S_ARBURST ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARBURST ),
        .FIC_1_AXI4_S_ARQOS   ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARQOS ),
        .FIC_1_AXI4_S_ARLOCK  ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLOCK ),
        .FIC_1_AXI4_S_ARCACHE ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARCACHE ),
        .FIC_1_AXI4_S_ARPROT  ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARPROT ),
        .FIC_1_AXI4_S_ARVALID ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARVALID ),
        .FIC_1_AXI4_S_RREADY  ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RREADY ),
        .FIC_2_ACLK           ( FIC_2_ACLK ),
        .FIC_2_AXI4_S_AWID    ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWID ),
        .FIC_2_AXI4_S_AWADDR  ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWADDR ),
        .FIC_2_AXI4_S_AWLEN   ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLEN ),
        .FIC_2_AXI4_S_AWSIZE  ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWSIZE ),
        .FIC_2_AXI4_S_AWBURST ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWBURST ),
        .FIC_2_AXI4_S_AWLOCK  ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLOCK ),
        .FIC_2_AXI4_S_AWCACHE ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWCACHE ),
        .FIC_2_AXI4_S_AWQOS   ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWQOS ),
        .FIC_2_AXI4_S_AWPROT  ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWPROT ),
        .FIC_2_AXI4_S_AWVALID ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWVALID ),
        .FIC_2_AXI4_S_WDATA   ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WDATA ),
        .FIC_2_AXI4_S_WSTRB   ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WSTRB ),
        .FIC_2_AXI4_S_WLAST   ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WLAST ),
        .FIC_2_AXI4_S_WVALID  ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WVALID ),
        .FIC_2_AXI4_S_BREADY  ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BREADY ),
        .FIC_2_AXI4_S_ARID    ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARID ),
        .FIC_2_AXI4_S_ARADDR  ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARADDR ),
        .FIC_2_AXI4_S_ARLEN   ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLEN ),
        .FIC_2_AXI4_S_ARSIZE  ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARSIZE ),
        .FIC_2_AXI4_S_ARBURST ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARBURST ),
        .FIC_2_AXI4_S_ARLOCK  ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLOCK ),
        .FIC_2_AXI4_S_ARCACHE ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARCACHE ),
        .FIC_2_AXI4_S_ARQOS   ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARQOS ),
        .FIC_2_AXI4_S_ARPROT  ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARPROT ),
        .FIC_2_AXI4_S_ARVALID ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARVALID ),
        .FIC_2_AXI4_S_RREADY  ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RREADY ),
        .FIC_3_PCLK           ( FIC_3_PCLK ),
        .FIC_3_APB_M_PRDATA   ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PRDATA ),
        .FIC_3_APB_M_PREADY   ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PREADY ),
        .FIC_3_APB_M_PSLVERR  ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PSLVERR ),
        .MMUART_1_DCD_F2M     ( VCC_net ),
        .MMUART_1_RI_F2M      ( VCC_net ),
        .MMUART_1_DSR_F2M     ( VCC_net ),
        .MMUART_1_CTS_F2M     ( M2_UART_CTS ),
        .MMUART_1_RXD_F2M     ( M2_UART_RXD ),
        .MMUART_2_RXD_F2M     ( MMUART_2_RXD ),
        .MMUART_3_RXD_F2M     ( MMUART_3_RXD ),
        .MMUART_4_RXD_F2M     ( MMUART_4_RXD ),
        .SPI_0_SS_F2M         ( GND_net ),
        .SPI_0_DI_F2M         ( SPI_0_DI ),
        .SPI_0_CLK_F2M        ( GND_net ),
        .SPI_1_SS_F2M         ( GND_net ),
        .SPI_1_DI_F2M         ( SPI_1_DI ),
        .SPI_1_CLK_F2M        ( GND_net ),
        .I2C_0_SCL_F2M        ( I2C0_SCL_BIBUF_Y ),
        .I2C_0_SDA_F2M        ( I2C0_SDA_BIBUF_Y ),
        .GPIO_2_F2M_31        ( SD_DET ),
        .GPIO_2_F2M_27        ( GPIO_2_F2M_slice_0 ),
        .GPIO_2_F2M_26        ( GPIO_2_F2M_slice_1 ),
        .GPIO_2_F2M_25        ( GPIO_2_F2M_slice_2 ),
        .GPIO_2_F2M_24        ( GPIO_2_F2M_slice_3 ),
        .GPIO_2_F2M_23        ( GPIO_2_F2M_slice_4 ),
        .GPIO_2_F2M_22        ( GPIO_2_F2M_slice_5 ),
        .GPIO_2_F2M_21        ( GPIO_2_F2M_slice_6 ),
        .GPIO_2_F2M_20        ( GPIO_2_F2M_slice_7 ),
        .GPIO_2_F2M_19        ( GPIO_2_F2M_slice_8 ),
        .GPIO_2_F2M_18        ( GPIO_2_F2M_slice_9 ),
        .GPIO_2_F2M_17        ( GPIO_2_F2M_slice_10 ),
        .GPIO_2_F2M_16        ( GPIO_2_F2M_slice_11 ),
        .GPIO_2_F2M_15        ( GPIO_2_F2M_slice_12 ),
        .GPIO_2_F2M_14        ( GPIO_2_F2M_slice_13 ),
        .GPIO_2_F2M_13        ( GPIO_2_F2M_slice_14 ),
        .GPIO_2_F2M_12        ( GPIO_2_F2M_slice_15 ),
        .GPIO_2_F2M_11        ( GPIO_2_F2M_slice_16 ),
        .GPIO_2_F2M_10        ( GPIO_2_F2M_slice_17 ),
        .GPIO_2_F2M_9         ( GPIO_2_F2M_slice_18 ),
        .GPIO_2_F2M_8         ( GPIO_2_F2M_slice_19 ),
        .GPIO_2_F2M_7         ( GPIO_2_F2M_slice_20 ),
        .GPIO_2_F2M_6         ( GPIO_2_F2M_slice_21 ),
        .GPIO_2_F2M_5         ( GPIO_2_F2M_slice_22 ),
        .GPIO_2_F2M_4         ( GPIO_2_F2M_slice_23 ),
        .GPIO_2_F2M_3         ( GPIO_2_F2M_slice_24 ),
        .GPIO_2_F2M_2         ( GPIO_2_F2M_slice_25 ),
        .GPIO_2_F2M_1         ( GPIO_2_F2M_slice_26 ),
        .GPIO_2_F2M_0         ( GPIO_2_F2M_slice_27 ),
        .MAC_1_MDI_F2M        ( MAC_1_MDI_F2M ),
        .MSS_INT_F2M          ( MSS_INT_F2M_net_0 ),
        .MSS_RESET_N_F2M      ( VCC_net ),
        .MMUART_0_RXD         ( UART0_RXD ),
        .GPIO_0_13_IN         ( USER_BUTTON ),
        .GPIO_1_20_IN         ( ADC_IRQn ),
        .GPIO_1_23_IN         ( USB_OCn ),
        .USB_CLK              ( USB_CLK ),
        .USB_DIR              ( USB_DIR ),
        .USB_NXT              ( USB_NXT ),
        .EMMC_STRB            ( EMMC_STRB ),
        .SGMII_RX1_P          ( SGMII_RX1_P ),
        .SGMII_RX1_N          ( SGMII_RX1_N ),
        .SGMII_RX0_P          ( SGMII_RX0_P ),
        .SGMII_RX0_N          ( SGMII_RX0_N ),
        .REFCLK               ( REFCLK ),
        .REFCLK_N             ( REFCLK_N ),
        // Outputs
        .FIC_0_DLL_LOCK_M2F   ( PF_SOC_MSS_FIC_0_DLL_LOCK_M2F ),
        .FIC_1_DLL_LOCK_M2F   ( PF_SOC_MSS_FIC_1_DLL_LOCK_M2F ),
        .FIC_2_DLL_LOCK_M2F   ( PF_SOC_MSS_FIC_2_DLL_LOCK_M2F ),
        .FIC_3_DLL_LOCK_M2F   ( PF_SOC_MSS_FIC_3_DLL_LOCK_M2F ),
        .FIC_0_AXI4_M_AWID    ( FIC_0_AXI4_INITIATOR_AWID ),
        .FIC_0_AXI4_M_AWADDR  ( FIC_0_AXI4_INITIATOR_AWADDR ),
        .FIC_0_AXI4_M_AWLEN   ( FIC_0_AXI4_INITIATOR_AWLEN ),
        .FIC_0_AXI4_M_AWSIZE  ( FIC_0_AXI4_INITIATOR_AWSIZE ),
        .FIC_0_AXI4_M_AWBURST ( FIC_0_AXI4_INITIATOR_AWBURST ),
        .FIC_0_AXI4_M_AWLOCK  ( FIC_0_AXI4_INITIATOR_AWLOCK ),
        .FIC_0_AXI4_M_AWQOS   ( FIC_0_AXI4_INITIATOR_AWQOS ),
        .FIC_0_AXI4_M_AWCACHE ( FIC_0_AXI4_INITIATOR_AWCACHE ),
        .FIC_0_AXI4_M_AWPROT  ( FIC_0_AXI4_INITIATOR_AWPROT ),
        .FIC_0_AXI4_M_AWVALID ( FIC_0_AXI4_INITIATOR_AWVALID ),
        .FIC_0_AXI4_M_WDATA   ( FIC_0_AXI4_INITIATOR_WDATA ),
        .FIC_0_AXI4_M_WSTRB   ( FIC_0_AXI4_INITIATOR_WSTRB ),
        .FIC_0_AXI4_M_WLAST   ( FIC_0_AXI4_INITIATOR_WLAST ),
        .FIC_0_AXI4_M_WVALID  ( FIC_0_AXI4_INITIATOR_WVALID ),
        .FIC_0_AXI4_M_BREADY  ( FIC_0_AXI4_INITIATOR_BREADY ),
        .FIC_0_AXI4_M_ARID    ( FIC_0_AXI4_INITIATOR_ARID ),
        .FIC_0_AXI4_M_ARADDR  ( FIC_0_AXI4_INITIATOR_ARADDR ),
        .FIC_0_AXI4_M_ARLEN   ( FIC_0_AXI4_INITIATOR_ARLEN ),
        .FIC_0_AXI4_M_ARSIZE  ( FIC_0_AXI4_INITIATOR_ARSIZE ),
        .FIC_0_AXI4_M_ARBURST ( FIC_0_AXI4_INITIATOR_ARBURST ),
        .FIC_0_AXI4_M_ARLOCK  ( FIC_0_AXI4_INITIATOR_ARLOCK ),
        .FIC_0_AXI4_M_ARQOS   ( FIC_0_AXI4_INITIATOR_ARQOS ),
        .FIC_0_AXI4_M_ARCACHE ( FIC_0_AXI4_INITIATOR_ARCACHE ),
        .FIC_0_AXI4_M_ARPROT  ( FIC_0_AXI4_INITIATOR_ARPROT ),
        .FIC_0_AXI4_M_ARVALID ( FIC_0_AXI4_INITIATOR_ARVALID ),
        .FIC_0_AXI4_M_RREADY  ( FIC_0_AXI4_INITIATOR_RREADY ),
        .FIC_0_AXI4_S_AWREADY ( FIC_0_AXI4_TARGET_AWREADY ),
        .FIC_0_AXI4_S_WREADY  ( FIC_0_AXI4_TARGET_WREADY ),
        .FIC_0_AXI4_S_BID     ( FIC_0_AXI4_TARGET_BID ),
        .FIC_0_AXI4_S_BRESP   ( FIC_0_AXI4_TARGET_BRESP ),
        .FIC_0_AXI4_S_BVALID  ( FIC_0_AXI4_TARGET_BVALID ),
        .FIC_0_AXI4_S_ARREADY ( FIC_0_AXI4_TARGET_ARREADY ),
        .FIC_0_AXI4_S_RID     ( FIC_0_AXI4_TARGET_RID ),
        .FIC_0_AXI4_S_RDATA   ( FIC_0_AXI4_TARGET_RDATA ),
        .FIC_0_AXI4_S_RRESP   ( FIC_0_AXI4_TARGET_RRESP ),
        .FIC_0_AXI4_S_RLAST   ( FIC_0_AXI4_TARGET_RLAST ),
        .FIC_0_AXI4_S_RVALID  ( FIC_0_AXI4_TARGET_RVALID ),
        .FIC_1_AXI4_M_AWID    ( FIC_1_AXI4_INITIATOR_AWID ),
        .FIC_1_AXI4_M_AWADDR  ( FIC_1_AXI4_INITIATOR_AWADDR ),
        .FIC_1_AXI4_M_AWLEN   ( FIC_1_AXI4_INITIATOR_AWLEN ),
        .FIC_1_AXI4_M_AWSIZE  ( FIC_1_AXI4_INITIATOR_AWSIZE ),
        .FIC_1_AXI4_M_AWBURST ( FIC_1_AXI4_INITIATOR_AWBURST ),
        .FIC_1_AXI4_M_AWLOCK  ( FIC_1_AXI4_INITIATOR_AWLOCK ),
        .FIC_1_AXI4_M_AWQOS   ( FIC_1_AXI4_INITIATOR_AWQOS ),
        .FIC_1_AXI4_M_AWCACHE ( FIC_1_AXI4_INITIATOR_AWCACHE ),
        .FIC_1_AXI4_M_AWPROT  ( FIC_1_AXI4_INITIATOR_AWPROT ),
        .FIC_1_AXI4_M_AWVALID ( FIC_1_AXI4_INITIATOR_AWVALID ),
        .FIC_1_AXI4_M_WDATA   ( FIC_1_AXI4_INITIATOR_WDATA ),
        .FIC_1_AXI4_M_WSTRB   ( FIC_1_AXI4_INITIATOR_WSTRB ),
        .FIC_1_AXI4_M_WLAST   ( FIC_1_AXI4_INITIATOR_WLAST ),
        .FIC_1_AXI4_M_WVALID  ( FIC_1_AXI4_INITIATOR_WVALID ),
        .FIC_1_AXI4_M_BREADY  ( FIC_1_AXI4_INITIATOR_BREADY ),
        .FIC_1_AXI4_M_ARID    ( FIC_1_AXI4_INITIATOR_ARID ),
        .FIC_1_AXI4_M_ARADDR  ( FIC_1_AXI4_INITIATOR_ARADDR ),
        .FIC_1_AXI4_M_ARLEN   ( FIC_1_AXI4_INITIATOR_ARLEN ),
        .FIC_1_AXI4_M_ARSIZE  ( FIC_1_AXI4_INITIATOR_ARSIZE ),
        .FIC_1_AXI4_M_ARBURST ( FIC_1_AXI4_INITIATOR_ARBURST ),
        .FIC_1_AXI4_M_ARLOCK  ( FIC_1_AXI4_INITIATOR_ARLOCK ),
        .FIC_1_AXI4_M_ARQOS   ( FIC_1_AXI4_INITIATOR_ARQOS ),
        .FIC_1_AXI4_M_ARCACHE ( FIC_1_AXI4_INITIATOR_ARCACHE ),
        .FIC_1_AXI4_M_ARPROT  ( FIC_1_AXI4_INITIATOR_ARPROT ),
        .FIC_1_AXI4_M_ARVALID ( FIC_1_AXI4_INITIATOR_ARVALID ),
        .FIC_1_AXI4_M_RREADY  ( FIC_1_AXI4_INITIATOR_RREADY ),
        .FIC_1_AXI4_S_AWREADY ( FIC_1_AXI4_TARGET_AWREADY ),
        .FIC_1_AXI4_S_WREADY  ( FIC_1_AXI4_TARGET_WREADY ),
        .FIC_1_AXI4_S_BID     ( FIC_1_AXI4_TARGET_BID ),
        .FIC_1_AXI4_S_BRESP   ( FIC_1_AXI4_TARGET_BRESP ),
        .FIC_1_AXI4_S_BVALID  ( FIC_1_AXI4_TARGET_BVALID ),
        .FIC_1_AXI4_S_ARREADY ( FIC_1_AXI4_TARGET_ARREADY ),
        .FIC_1_AXI4_S_RID     ( FIC_1_AXI4_TARGET_RID ),
        .FIC_1_AXI4_S_RDATA   ( FIC_1_AXI4_TARGET_RDATA ),
        .FIC_1_AXI4_S_RRESP   ( FIC_1_AXI4_TARGET_RRESP ),
        .FIC_1_AXI4_S_RLAST   ( FIC_1_AXI4_TARGET_RLAST ),
        .FIC_1_AXI4_S_RVALID  ( FIC_1_AXI4_TARGET_RVALID ),
        .FIC_2_AXI4_S_AWREADY ( FIC_2_AXI4_TARGET_AWREADY ),
        .FIC_2_AXI4_S_WREADY  ( FIC_2_AXI4_TARGET_WREADY ),
        .FIC_2_AXI4_S_BID     ( FIC_2_AXI4_TARGET_BID ),
        .FIC_2_AXI4_S_BRESP   ( FIC_2_AXI4_TARGET_BRESP ),
        .FIC_2_AXI4_S_BVALID  ( FIC_2_AXI4_TARGET_BVALID ),
        .FIC_2_AXI4_S_ARREADY ( FIC_2_AXI4_TARGET_ARREADY ),
        .FIC_2_AXI4_S_RID     ( FIC_2_AXI4_TARGET_RID ),
        .FIC_2_AXI4_S_RDATA   ( FIC_2_AXI4_TARGET_RDATA ),
        .FIC_2_AXI4_S_RRESP   ( FIC_2_AXI4_TARGET_RRESP ),
        .FIC_2_AXI4_S_RLAST   ( FIC_2_AXI4_TARGET_RLAST ),
        .FIC_2_AXI4_S_RVALID  ( FIC_2_AXI4_TARGET_RVALID ),
        .FIC_3_APB_M_PSEL     ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PSELx ),
        .FIC_3_APB_M_PADDR    ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PADDR ),
        .FIC_3_APB_M_PWRITE   ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PWRITE ),
        .FIC_3_APB_M_PENABLE  ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PENABLE ),
        .FIC_3_APB_M_PSTRB    ( FIC_3_APB_M_PSTRB_net_0 ),
        .FIC_3_APB_M_PWDATA   ( PF_SOC_MSS_FIC_3_APB_INITIATOR_PWDATA ),
        .MMUART_1_DTR_M2F     (  ),
        .MMUART_1_RTS_M2F     ( M2_UART_RTS_net_0 ),
        .MMUART_1_TXD_M2F     ( M2_UART_TXD_net_0 ),
        .MMUART_1_TXD_OE_M2F  (  ),
        .MMUART_2_TXD_M2F     ( MMUART_2_TXD_net_0 ),
        .MMUART_3_TXD_M2F     ( MMUART_3_TXD_net_0 ),
        .MMUART_4_TXD_M2F     ( MMUART_4_TXD_net_0 ),
        .SPI_0_SS1_M2F        ( SPI_0_SS1_net_0 ),
        .SPI_0_SS1_OE_M2F     (  ),
        .SPI_1_SS1_M2F        ( SPI_1_SS1_net_0 ),
        .SPI_1_SS1_OE_M2F     (  ),
        .SPI_0_DO_M2F         ( SPI_0_DO_net_0 ),
        .SPI_0_DO_OE_M2F      (  ),
        .SPI_0_CLK_M2F        ( SPI_0_CLK_net_0 ),
        .SPI_0_CLK_OE_M2F     (  ),
        .SPI_1_DO_M2F         ( SPI_1_DO_net_0 ),
        .SPI_1_DO_OE_M2F      (  ),
        .SPI_1_CLK_M2F        ( SPI_1_CLK_net_0 ),
        .SPI_1_CLK_OE_M2F     (  ),
        .I2C_0_SCL_OE_M2F     ( PF_SOC_MSS_I2C_0_SCL_OE_M2F ),
        .I2C_0_SDA_OE_M2F     ( PF_SOC_MSS_I2C_0_SDA_OE_M2F ),
        .GPIO_2_M2F_30        ( VIO_ENABLE_net_0 ),
        .GPIO_2_M2F_29        ( M2_W_DISABLE2_net_0 ),
        .GPIO_2_M2F_28        ( M2_W_DISABLE1_net_0 ),
        .GPIO_2_M2F_27        ( GPIO_2_M2F_net_0 ),
        .GPIO_2_M2F_26        ( GPIO_2_M2F_0 ),
        .GPIO_2_M2F_25        ( GPIO_2_M2F_1 ),
        .GPIO_2_M2F_24        ( GPIO_2_M2F_2 ),
        .GPIO_2_M2F_23        ( GPIO_2_M2F_3 ),
        .GPIO_2_M2F_22        ( GPIO_2_M2F_4 ),
        .GPIO_2_M2F_21        ( GPIO_2_M2F_5 ),
        .GPIO_2_M2F_20        ( GPIO_2_M2F_6 ),
        .GPIO_2_M2F_19        ( GPIO_2_M2F_7 ),
        .GPIO_2_M2F_18        ( GPIO_2_M2F_8 ),
        .GPIO_2_M2F_17        ( GPIO_2_M2F_9 ),
        .GPIO_2_M2F_16        ( GPIO_2_M2F_10 ),
        .GPIO_2_M2F_15        ( GPIO_2_M2F_11 ),
        .GPIO_2_M2F_14        ( GPIO_2_M2F_12 ),
        .GPIO_2_M2F_13        ( GPIO_2_M2F_13 ),
        .GPIO_2_M2F_12        ( GPIO_2_M2F_14 ),
        .GPIO_2_M2F_11        ( GPIO_2_M2F_15 ),
        .GPIO_2_M2F_10        ( GPIO_2_M2F_16 ),
        .GPIO_2_M2F_9         ( GPIO_2_M2F_17 ),
        .GPIO_2_M2F_8         ( GPIO_2_M2F_18 ),
        .GPIO_2_M2F_7         ( GPIO_2_M2F_19 ),
        .GPIO_2_M2F_6         ( GPIO_2_M2F_20 ),
        .GPIO_2_M2F_5         ( GPIO_2_M2F_21 ),
        .GPIO_2_M2F_4         ( GPIO_2_M2F_22 ),
        .GPIO_2_M2F_3         ( GPIO_2_M2F_23 ),
        .GPIO_2_M2F_2         ( GPIO_2_M2F_24 ),
        .GPIO_2_M2F_1         ( GPIO_2_M2F_25 ),
        .GPIO_2_M2F_0         ( GPIO_2_M2F_26 ),
        .GPIO_2_OE_M2F_27     ( GPIO_2_OE_M2F_net_0 ),
        .GPIO_2_OE_M2F_26     ( GPIO_2_OE_M2F_0 ),
        .GPIO_2_OE_M2F_25     ( GPIO_2_OE_M2F_1 ),
        .GPIO_2_OE_M2F_24     ( GPIO_2_OE_M2F_2 ),
        .GPIO_2_OE_M2F_23     ( GPIO_2_OE_M2F_3 ),
        .GPIO_2_OE_M2F_22     ( GPIO_2_OE_M2F_4 ),
        .GPIO_2_OE_M2F_21     ( GPIO_2_OE_M2F_5 ),
        .GPIO_2_OE_M2F_20     ( GPIO_2_OE_M2F_6 ),
        .GPIO_2_OE_M2F_19     ( GPIO_2_OE_M2F_7 ),
        .GPIO_2_OE_M2F_18     ( GPIO_2_OE_M2F_8 ),
        .GPIO_2_OE_M2F_17     ( GPIO_2_OE_M2F_9 ),
        .GPIO_2_OE_M2F_16     ( GPIO_2_OE_M2F_10 ),
        .GPIO_2_OE_M2F_15     ( GPIO_2_OE_M2F_11 ),
        .GPIO_2_OE_M2F_14     ( GPIO_2_OE_M2F_12 ),
        .GPIO_2_OE_M2F_13     ( GPIO_2_OE_M2F_13 ),
        .GPIO_2_OE_M2F_12     ( GPIO_2_OE_M2F_14 ),
        .GPIO_2_OE_M2F_11     ( GPIO_2_OE_M2F_15 ),
        .GPIO_2_OE_M2F_10     ( GPIO_2_OE_M2F_16 ),
        .GPIO_2_OE_M2F_9      ( GPIO_2_OE_M2F_17 ),
        .GPIO_2_OE_M2F_8      ( GPIO_2_OE_M2F_18 ),
        .GPIO_2_OE_M2F_7      ( GPIO_2_OE_M2F_19 ),
        .GPIO_2_OE_M2F_6      ( GPIO_2_OE_M2F_20 ),
        .GPIO_2_OE_M2F_5      ( GPIO_2_OE_M2F_21 ),
        .GPIO_2_OE_M2F_4      ( GPIO_2_OE_M2F_22 ),
        .GPIO_2_OE_M2F_3      ( GPIO_2_OE_M2F_23 ),
        .GPIO_2_OE_M2F_2      ( GPIO_2_OE_M2F_24 ),
        .GPIO_2_OE_M2F_1      ( GPIO_2_OE_M2F_25 ),
        .GPIO_2_OE_M2F_0      ( GPIO_2_OE_M2F_26 ),
        .MAC_1_MDO_M2F        ( MAC_1_MDO_M2F_net_0 ),
        .MAC_1_MDO_OE_M2F     ( MAC_1_MDO_OE_M2F_net_0 ),
        .MAC_1_MDC_M2F        ( MAC_1_MDC_M2F_net_0 ),
        .MSS_INT_M2F          (  ),
        .PLL_CPU_LOCK_M2F     (  ),
        .PLL_DDR_LOCK_M2F     (  ),
        .PLL_SGMII_LOCK_M2F   (  ),
        .MSS_RESET_N_M2F      ( MSS_RESET_N_M2F_net_0 ),
        .MMUART_0_TXD         ( UART0_TXD_net_0 ),
        .MAC_0_MDC            ( PHY_MDC_net_0 ),
        .GPIO_0_12_OUT        ( SD_CARD_CS_net_0 ),
        .USB_STP              ( USB_STP_net_0 ),
        .QSPI_SS0             ( ADC_CSn_net_0 ),
        .QSPI_CLK             ( ADC_SCK_net_0 ),
        .EMMC_CLK             ( EMMC_CLK_net_0 ),
        .EMMC_RSTN            ( EMMC_RSTN_net_0 ),
        .SGMII_TX1_P          ( SGMII_TX1_P_net_0 ),
        .SGMII_TX1_N          ( SGMII_TX1_N_net_0 ),
        .SGMII_TX0_P          ( SGMII_TX0_P_net_0 ),
        .SGMII_TX0_N          ( SGMII_TX0_N_net_0 ),
        .DM                   ( DM_net_0 ),
        .RESET_N              ( RESET_N_net_0 ),
        .ODT                  ( ODT_net_0 ),
        .CKE                  ( CKE_net_0 ),
        .CS                   ( CS_net_0 ),
        .CK                   ( CK_net_0 ),
        .CK_N                 ( CK_N_net_0 ),
        .CA                   ( CA_net_0 ),
        // Inouts
        .I2C_1_SCL            ( I2C_1_SCL ),
        .I2C_1_SDA            ( I2C_1_SDA ),
        .MAC_0_MDIO           ( PHY_MDIO ),
        .USB_DATA0            ( USB_DATA0 ),
        .USB_DATA1            ( USB_DATA1 ),
        .USB_DATA2            ( USB_DATA2 ),
        .USB_DATA3            ( USB_DATA3 ),
        .USB_DATA4            ( USB_DATA4 ),
        .USB_DATA5            ( USB_DATA5 ),
        .USB_DATA6            ( USB_DATA6 ),
        .USB_DATA7            ( USB_DATA7 ),
        .QSPI_DATA0           ( ADC_MOSI ),
        .QSPI_DATA1           ( ADC_MISO ),
        .EMMC_CMD             ( EMMC_CMD ),
        .EMMC_DATA0           ( EMMC_DATA0 ),
        .EMMC_DATA1           ( EMMC_DATA1 ),
        .EMMC_DATA2           ( EMMC_DATA2 ),
        .EMMC_DATA3           ( EMMC_DATA3 ),
        .EMMC_DATA4           ( EMMC_DATA4 ),
        .EMMC_DATA5           ( EMMC_DATA5 ),
        .EMMC_DATA6           ( EMMC_DATA6 ),
        .EMMC_DATA7           ( EMMC_DATA7 ),
        .DQ                   ( DQ ),
        .DQS                  ( DQS ),
        .DQS_N                ( DQS_N ) 
        );


endmodule
